��   ��A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����DCSS_C�PC_T  �4 $COMM�ENT $�ENABLE � $MODJG�RP_NUMKL�\  $U�FRM\] _VT�X M �   �$Y�Z1K �$Z2�STOP�_TYPKDSB�IO�IDXKE�NBL_CALM�D�USE_PR�EDIC? �EL�AY_TIMJS�PEED_CTR�LKOVR_LI�M? p D� L�0��UTOOi��O^*+&S. � 8J\TC�u
!���p\� E&|Y0  � �CHG_SIZ�O$AP!�E�DIS�]$!�!C_+{#s%O#J�p 	]$Jd#� �&s"�"�{#�)�$�'�_SE�EXPAN#N��  ,$STAT�/ DFP_�BASE 5$0K$4!� .6�_V7>H73��&J>- � }�n\AXS\UP��LW�7������d4r � < w?�?�?��?�?��//	0&ELE}M/ T �&B.2NO�G]@%CN�HA�DF#� $DATA)a6e0 � PJ�@ �2 
&P5� �� 1U*n   _VSiSZbRj0RjR(�VyT(�R%S�{TROBOT�X�SARo�U�V$C�UR_��R DSE�TU4"	 �bAI�SP_MGN�I?NP_ASSe#� PB!� `CiH�77`e��.fXc1�CONFIG_CHK`E�_PO* }dSHR�ST�gM^#/eOT�HERRBT�j_G]�R�dTv �ku,�chT1r
0R HpLH�d� 0  lt<xNe'AVRFYhH�^t�5�1� ��W��_A$R�4S;PH/ (G%�Q�Q�Q3wB;OX/ 8�@F!��F!�G �r{�zT�UIRi@  �,�F�pER%@2� $�p -L�_SF��D(��ZN/ 0 �IF(@�p��Z_��0�_�0wu0 � @�Q7yv	
�� _�$$CL` �2�����Q��Q��V�ERSION���  �Z��$' 2 �Q�  C�ell Box �In��*�h� ���m�����E�"� œ�����E� ŷ�����?Ĩ� D�ğ�����  d����Cz  ����:����JackpotT�Out_�q�w�,�����c��@���?�^� DH��Κ�@ȯ+���9�'��I�Incomi�ng[�n�����a � E	����D\ G �ȩ���ޡ�ÿ -���;�)�G�H�l� {���oϬ�������h����%�7�I�MiddleT�h�~���?9  �8`L߫�?C�&få��Οl�
��`15���C��1�G�Left Side�`�u��ߐ�O;� E�߭�CԐ�����Д�  D���������D�B�>D�Righg�z� �������ྱ���� ��Q��%�K�9O��ICK SLOW�DOW�z�߃�"ؐ�������ě����n�0BW�b�d�J2 SlowdowZ�������������[�C ې����1/E/_�h�z����D�����/ #/5/?I?Sπ?wω� ���?�?�?�??1? C?U?g?|O�O�?�?�O �?�O�O�OO-O?OQO�f_Y�pick d?cs tesb��)d����_��Ö@P�P�_`��ې�Qo_ ._@_R_TorO�o�O�O �O�o�o�o	o*o<o No`oro���o�o� �o���&8J\ ������p��̏ ��"�4�F�l�j�|� �����ďٟ���� �0�B�T�f�{����� ����������,� >�P�v�d��������� ί����(�:�L� ^�p��ϔ��ϸ�ʿ�� ���'�6�H�Z� � nߐϥߴ��������� �#�2�D�V�h�zߏ� �߳����������� 1�@�R�d�v�x���� ���������-<� N�`�r��������� ���)�J\ n�;����� ��%/7/FXj� ���/@/���// !?3?B/T/f/x/�/�? �/�?�/�/�??	O/O AOP?b?t?�?�O�?�O �?�?�?_O+_=_LO ^OpO�O�O�_�O�_�O �Oo_'o9oKoZ_l_ ~_$o�o�_�o�_�_�_  o5GVohozo�o �o��o��o�o� 1�C�U�dv���� �ӏ��*��
�?��Q�`�r�����������$DCSS_CS�C 2��ۑ�Q  P�100% S�afe Spee�}�b�l�F@
�,�ł�j�di1��j�C���'�,�
����i�����d�����ԯ 5���Y��i���R��� v�׿��������1� U��y�<ϝ�`��τ� ���Ϻ����?��c� &߇�J�\߽߀��ߤ� ���)���9�_�"���F��j����ΔGR�P 2ۛ ��ÄC��\En�њC  E5�� 	��5�ǀ#� \�G���k��������� ������F1j U�y����� �0T?xc ������/� />/)/b/M/�/�/�/ u/�/�/�/�/?(?? L?7?p?�?�?_?�?�? �?�? O�?�?6O!OZO lO~OIO�O�O�O�O�O �O_ __D_V_h_3_ �_w_�_�_�_�_�_�_��_.oŝGSTAT� 2ۙ-��<� ��?]����  G9�E�����f�]�9����;���;˒j��1�D�J�O��ODI�ۑ`<jf��9��
{�2�%DN4�t?׀  �a��`4���ZC��?��� Ɓۑje����+<��?t��S�tg�<��� ���e�i���y�>E��D��Y{�i>Hw�����?}�s<��	f�a�����}��<��=�>X�A�0���9��D�9_�{b�+��?�}�Bt�Jq�� ���,�����D�.�U�kD~�6�i?����;�~-�=p�p,;�ϫ������ː?�b�no�o �o�gە�0�ە�\� n�H��������j�`i ҏk�z����	�+� -�?�a���u���ş�� ��ߟះ�=�O���[� ��_�q���ͯÏ��� %��-��%�G�u�[� }��������ǿٿ�� )�+�ѯkϝ�Wϡϳ����������?]�����`9�R���6�p����3 ;��K;����p0�`k�O?��DI��o�a���cB�g���k����k�<����`}�th�<��򾗘Vnf���2p� p��{F�p�2p��<��:t�}��<���>�V�A�?Q�9뎏Vpv{u��+�=np/���~��ѽ �	�s� ��pU�U�D~��4�|�A�;~��=�s�������˓��p1�(�
��.��� �������������8� J��2�t�Fό����� ����������(@ ^DVx�L��� ��0
Tf\� �������� /�/D/*/</^/�/ r/�/�/�/n?6�/ :?L?&?p?�?\?z�� 2�D�V�h�zߌߞ߰� ��������
��.�@� R��O�?�?�?d?V_h_ ^?t_�_x_�_�_�_� �/o�/(oFo,o>o`o �oto�o�o�o�o�o�o �oB�/r��_p ������_F,� Z$�F�t�Z�|����� ����Ə؏��(��0� ^�D�
������֟� ����_(_�?�? �?OO(O:OLO^OpO �O�O�O�O�O�O�O`� B�T�f� ������ :��&�pς��j��� ~�����������*�� 2�`�F�xߖ�|ߎ߰� �߄�� �R��V�h� B������������ ������F�,�N�|� b�t������������� ��<n�(r�^� ����Ŀj�|����� ��į֯�����0� B�T�f�x������ ��/�/��/�/�/ �/??��H?`? ~?d?v?�?�?�?�?�? �?O2OO*OLOzO  �O�O�/�O�O_�O(_ :_0?~Od_�O\_~_�_ �_�_�_�_�_o�_o 2o`oFoho�o|oB_�o 
_�o �oDV0 N/`/*<N` r������� //&/��z��8 *�<�2H�r�L�^��� ��T_�o䟶o��� � �4�b�H�j���~��� ί��Ư���oF�X� ��D�����z�Ŀֿ̟ � �.����H�.�P� ~�dφϴϚϬ����� ���2��޿tߦ�`� �߼ߖ���������� ������� � 2�D�V�h�z������� 4��(�:������� ��������DV� >߀Rߘ���� ��4LjP b��X���&� */<//`/r/h��/ ��/�/�/�/�/? ? "?P?6?H?j?�?~?�? �?�?z/OB/�?FOXO 2O|O�OhO����>�P� b�t��������� ����(�:�L�^��_ �O�O�OpObotojO�o �o�o�o�o�o�/�? �?4R8Jl�� ������� � N��?~����o|�Ə؏ �����R�8�f�0� R���f���������� ҟ��4��<�j�P� ���ޏ�����ί��*�8��$DCSS_JPC 2"��Q ( �DRight� Side Cl�ear����C9�  @@��
#P>"QLefn��J�����Õ�����In j��������C*�� �����򰮶����!��/"�!R}�D�Ǝ��At Pic�k���A  ����$�
RH Jackpot��̕��C!���L�߇�� a�ݳkό�Sߡ��Ⱦ�Home J1���˿ٙ���f�f4���2��������������3��������#�3_�G���4a��K�P�����5����¤  ¤�����6������>���at �EOAT chg� ���B�ffB��R�f��/�@Fff@����_�~s��������(�������vߨ�t����b j��d���+�?�B�  B��bdsblB�� f����� �������2������$.�3J�
�'�"{4���"Q�s���5 a��� �j��6��� �B�>/�ߥ/�߮�~F�2 limiO�V.�B�
�P���# ��/�/?#P�/m? �/�?`?�?�?�?�?�? �?�?3OOAO&O{OJO �OnO�O�O�O�O_�O �OA__"_4_�_X_�_�|_�_�_�_J�SS��W�L  afe? Speed�_»Bȉ�H�1aG�a2&`to�o7�A8�� aaai��ro�o�_�ofa �o�o?c*� N�r����� �;�M��q�8���\� ����ݏ���ȏ%�� 3��m�4�F�X�j�ǟ ��럲��֟3���W� �{�B���f�x���� ������A��e�,� ��P���t�ѿ��߿�� �����s�:ϗ� ^ϻς��Ϧ����'� ��K��$�6ߓߥ�l� �ߐ��ߴ����5��� Y� �}�D��h���� ��������C�
�g� .���R���v������� ������?Qu< �`����� )�7q8J\�n����dMO�DEL 2k�x^!��$<��c�X B���fÈ  A`�  CHp �� ��o$F/X/�	p xp$6  ë$�/�/j&�t(� �/�/�&�!�%�#�9�!�hM7 b?9?K?�?o?�?�?�? �?�?O�?�?LO#O5O<GO�WJ3 �O=-M=C\�(s �s 3��� �@CW�CbO tO�O\O__e_<_N_ �_r_�_�_�_�_�_o �_oOo&o8oWo\ono`�o�o�o�o� �L�o�o\�oEWi {������� ��/�A���e�w�ď ������я���B�� +�x�%S�e�ҟM� ��͟���P�'�9� ��]�o���ί����� ۯ�:��#�5���Y� k������������ ۿ�ÿ1�Cϐ�g�y� �ϝϯ���������D� �-�z�Q�c�u߇ߙ� ��������.���)� ����#�Q�c�9��� �����<��%�7�I� [�m������������� ����!nEW� {��u������ F/|Se�� �����0/// f/=/O/a/�/�/�/�/ �/�/?�/??�t? =?O?�?�?�?�?�? �?�?�?O#OpOGOYO �O}O�O�O�O�O�O$_ �O_Z_1_C_U_g_y_ �_a?�_�?�_�_2o	o oho?oQocouo�o�o �o�o�o�o) ;M�q���� �����_`��_)� ;������ޏ��Ǐُ &����\�3�E���i� {���ڟ��ß���� F��/�A���e�w�M� _�q���������� +�=�O���s���ҿ�� ��Ϳ߿��P�'�9� ��]�oρϓϥϷ�� ����:�կ��'ߔ� �}ߏߡ߳������ ��H��1�C�U�g�y� ������������	� �-�z�Q�c���K�]� ����
����R) ;�_q���� ��<%rI [m������ &/������/%/�i/ {/�/�/�/�/�/�/�/ ??/?|?S?e?�?�? �?�?�?�?�?0OOO fO=OOOaO7/�O[/�O �OqO�O�O>__'_t_ K_]_o_�_�_�_�_�_ �_(o�_o#o5oGoYo �o}o�o�o�o�o�o�O 6�O�o~Ug� ������2�	� �h�?�Q���u����� 揽�Ϗ���R�)��;�M�f��$DCS�S_PSTAT �������Q   t�佐ɐПԐ  �Ν (t���x�����ʝ���ԟ;�� W�  t���k�損�����e�����¯p���鮦��SETUP 	��B�x�k��� 4���U�D�y�h�����T1SC 2
�f�m�Czk�ݿ�|ͺ�CP RȼD�D.L�^�  �ϔϦ�u������Ͻ� �$�6��Z�l�;�}� �ߴ߃��������� � 2�D��h�z��[�� �������
���.�@� R�!�v�����i����� ������<N` h�8ύ�&��� �/�Sew F������� /+/=//a/s/�/T/ �/�/�/�/�/?�/�/ 9?K??o?�?�?b?�? �?�?�?�?O#O�?GO YO(O}O�O�Op�O�O �OpO__1_ _U_g_ y_H_�_�_~_�_�_�_ �_o-o?oocouo�o Vo�o�o�o�o�o�o );Mq��d �������� I�[�*������r�Ǐ ُ돺O�!�3���W� i�{�J�������՟� ��ȟ�/�A��e�w� ��X������������ ֯+�=�O��s����� f���Ϳ߿����� 9�K�]�,ρϓϥ�t� �����ϼ��#�5�� Y�k���Lߡ߳߂��� �������1�C��g� y��Z��������� 	���-�?�Q� �u��� ��h��������� ��;M_.��� v����%� I[m<ߑ��< ����!/3/E// i/{/J/\/�/�/�/�/ �/?�//?A?S?"?w? �?�?j?�?�?�?�?O O�?=OOOaO0O�O�O �OxO�O�O�O�O_'_ �OK_]_o_>_�_�_�_ ��_�_�_�_#o5oGo oko}oLo�o�o�o�o �o�o�o1CU$ y�Zl���� 	���?�Q�c�2��� ����z�ϏᏰ��� )���M�_�q�@����� ����ݟ���_%�7� ���m��N�����ǯ ������ޯ3�E�W� &�{���\���ÿտ�� �����A�S�e�4� �ϛ�j�|����ϲ�� �+���O�a�s�Bߗ� �߻ߊ��������'��9���$DCSS�_TCPMAP � ���g��Q @ *����w�U����U	�
�������  U����U������������ �!��"�#�$�%��&�'�(�)��*�+�,�-��.�/�0�1��2�3�4�5��6�7�8�9��:�;�<�=��>�?�@W�U�IRO 2g��x�������� ������ 2DV hz�����������3EW i{������ �////A/S/e/� �/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?|/O�/ 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_�Y_k_}_O�_S�UI�ZN 2g�	 �x�v��_�_o� �_4oFoXoo|o�o�o oo�o�o�o�o0 �oTfx;��� ������>�P� �t�������m�Ώ�� ����(�:���^�p� ��Q�����ʟ��� � ��6�H�Z��/������q�Ưدꯩ_Z�U�FRM Rf����8�@�R��v� ��c����������Ͽ �*��N�`�;τϖ� qϺ��ϧ�����+� 8�J���n߀�[ߤ߶� ���������"���F� X�3�i���{����� �����#�0�B���f� x�S������������� ��,Pb=� �s����� (:�^pK�� �����/$/� H/Z/5/~/�/k/�/�/ �/�/�/
?2?D?? h?z?U?�?�?�?�?�? �?
OO�?@ORO-OvO �OcO�O�O�O�O�O? ?*_<_�O`_r_M_�_ �_�_�_�_�_oo�_ 8oJo%ono�o[o�o�o �o�o�o�o_"4�o XjE��{�� �����B�T�/� x���e���������� �,�ˏP�b�=��� ��s���Ο������ �:�L�'�p���]��� ����ܯ�ȧ