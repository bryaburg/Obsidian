��   !��A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETGX��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S�ETHOST� � �DNSS*� 8�D�FAC�E_NUM? $�DBG_LEVE�L�OM_NAM� !�* �D $PRIM�AR_IG !$?ALTERN1��<WAIT_TI�A �� FT�� @� LOG_�8	�CMO>$DNLD_FI:��SUBDIRCAP�����8 .� 4� H�A�DDRTYP�H NGTH��Y�z +LS�&$ROBOT2�PEER2� MA�SK4MRU~O�MGDEV��P�INFO� �$$$X �R�CMT A�$| ��QSIZ�X�� TATU�SWMAILSE�RV $PLA�N� <$LIN><$CLU����<$TO�P$C�C�&FR�&�JE�C�!�%ENB �� ALAR�!BF�TP�/3�V8 }S��$VAR79�M ON,6��,6A7PPL,6PA� -5�B +7POR��#_|12ALERT�&��2URL }>�3ATTAC��0�ERR_THRO��3US�9�!�8R0CqH- YDMAXN�S_�1�1AMOD�2AI� o 2A�� (1APWD � � LA �0�N�D)ATRYsFDE�LA�C2@�'`AERcSI�1A�'RO�ICLK�HMt0�'� �XML+ \3SGF�RM�3T� XOU̩3Z G_��COP c1V�3Q�'C�2-5R_AU�� � XR�N1oUPDXPC�OU�!SFO ?2 
$V~Wo��@YACC�H�QS�NAE$UMMY1Z�W2v$DM*	T �$DIS��S�MB�
 T &�	BCl@DCI2�AI&P6EXP9S�!�PAR� `�RANe@  ���QCL� �<(C�0�SPT9M
U� PWR�-h�CfSMo !l5��!�"%�7YD�P�% 0�fR�0z�eP� _DLV�$De\aNo3 
j��hX_!`�#Z_I�NDE,C_pOFF,� ~URnyD�*s��   t 9�!pMON��s�D��rHOU�#E�yA�v�q�v�q�vLOsCA� Y$N�0oH_HE��P�I"/  d	`A�RP�&�1F�W�_~ �I!Fap;F�A�D�01#�HO_Ȅ �R�2P$`�S�T;EL	% P K � !�0WO�` k�QE� LVt�k�2H#ICE��ڀ!� �$d� ? �������%
��
��`S$Q���  ��Z�$'0 �
�
��F����"�S�L�w�$� 24�T"�����e��� �4����ȟ����-�4�Ɵ��8�I�L����p_V`4�� S�z�������¯ԯ毀��
��.�@��� _?FLTR  �?�W �������!�ޛnx4�2ޛ8�{SHE`D 14�E P'��I�ٿ ��:���^�!ς�E� ��iϷ��ϟ� ���$� ��H��l�/�Aߢ�e� �߉��߭������D� �h�+��O��s�� ����
���.���R�� ^�9�����o������� ����<��r5 �Y�}��� �8�\�Cy�������PP�P_L�A1e�x/!1.9"0/��8%1I/�2551.�%@/��Q�7#2>/P.� d/v/�/�/�&3�/P.-0�/�/ ??�&4.?P.�0T?f?x?�?�&5�?P.@�?�?�?O�&6OP.�@�DOVOhOzOT�aP���t(�{��Ӱ��� OQ� ��N<0_ e_w_J_�_�_�_�_�_�_�P�_%o7oIoo moo�o�obo�o�o�o��N�o�T�5 |�
ZDT Status�oD�����}iRCon�nect: ir�c�t//alertb~���+��wt�Y�k�}��������2A�d�RJ������  ��$�6�H�Z�l�~��������ƟQs$$c�962b37a-�1ac0-eb2�a-f1c7-8�c6eb571d?066  (H��@l=�O�a�s���A
��X�'R��)z��`P��*s,P!T,$4� 񯨰*!߯��@�'� M�v�]�������п�� ��ۿ����N�5�r�4Y�����&%P7DM_Q	&+"?SMB 
&%U��#l��O���� �I��pb2����_CLNT �2&)9�4+t 	�|�#|j߯ߎߠ��� ��������Q�0�u�f������
.S�MTP_CTRL' R� P%��4� 	t��"�c���R���v�H��#|��N�Q�����7������ ��USTOM' ���&P� �TTCPIP����'xU"R�i EL$&%#Q�> H!TP	���rj3_tp�т��+ ��!K�CL�������!CRT.uR��!CONS�v�
�ib_s'mon~r