��   ��A��*SYST�EM*��V9.1�0170 9/�18/2019 A 	  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41�� d =RO &J_�  4 $:(F3IDX���_ICI  ��MIX_BG-<y
_NAMc gMODc_USd~�IFY_TI�� �MKR-�  $LIN�c   "_S�IZ��� �. �X $USE_FLC 3!�:&iF*SIMA7#Q�C#QBn'SCAN��AX�+IN�*I���_COUNrR�O( ��!_TMR�_VA�g# h>�ia �'` ����1�+WAR��$�H�!�#Nf3CH�PE�$,O�!PR�'Ioq6��OoATH-� P $ENA#BL+�0B�Tm��$$C�LASS  �����1��5��5��0VERS��7�  �Z��6/ �55�������@MF!�0�1RE��%�1{O��wO�O����#EI2.K!�O_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_oo�O+ �W?H9@ ���\j�0lo~o�i�ܧ � 2.I  4%BG���o���aP�|H%�o�g_A�oA  ewV���� �����=��.�@�c$"+ �kdK@����RA��X�� �1@fNʏ܏� �� $�6�H�Z�l�~����� ��RF_A��_A֟��� ��0�B�T�f�x���@�������4JM4��c6C!2�l��� /�A�S�e�w������� ��ѿ������(�:� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~ߐߢߴ������� ����2�D�V�h�z� ������������
� �'�@�R�d�v����� ����������#� <N`r���� ���&1J \n������ ��/"/-?X/j/ |/�/�/�/�/�/�/�/ ??0?3h�4�0v�g? @