��  Ij�A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����SBR_T �  | 	$S�VMTR_ID � $ROBO�T9$GRP�_NUM<AXIaSQ6K 6NFF�3 _PARAM�F	$�  �,$MD SPD�_LIT  &2j*� � �����$$CLASS  ���������� VER�SION��  �Z�$�'  1 � �T���R-�2000iC/1�25L���  �aiSR22/�4' 80A���
H1 DSP1�-S1��	P0�1.009,  	�  ���   ���# ������������
=��r�9  :�!a������ @H+ � ����� Y��� �v# < �����  �����&  �2�&���>A���$j���
"�����&��� �) 	���� ����������ߗ� ��A�����y���{����B� U K ���� �5� :?�����'b�
��E/�/�/�/�/��c�?��3?�C?U?g?��37X���=�����J���4]��<���\��cx�T�p?�?����0B30/3L2^2fx�ߜ���������~��%�����8 l�� ^߈�@����� ��*�*�����c	v� 5F����;�����Y�|���+�\, & �_��� �8$P�?�������\'w%��R��r(��c9	`�D 0��� ����#p�"=@��x��Ou_0�_�_�_3��_ ?0�_�_o��Z����5Y
��@��p����
��8m� �8u�����p��Toso�4�$�?0�?T3^�R"O4OFK��bZOlO~G����H��4��4��K|4D	 =���,����o(+�  , " �Bu|�O�����\'�
��h�q��-r(�6_H_Z_#�5�G�Y��-|h��_�� ��ŏ o�����1�l�o�o B10J�4Q4^4�o�m�:����(�����2�`8�	��� 0�� ��������yF�''@nq��`#�5���-�p_��� l8$�E���s���X���1��E	t�Ì�@��5P�!f� <�#S ��u�#'  �
�֯�����b	0�D;���fF� k�}�������ſ׿�LD�V� j�T5^15��������Ɵ؟��x��'�������������+ ��\�O`:"��Dn���[X}����R
�o�e✥�����ʯ�ߥ߷����-
(��H���#�5�G�Y��k�}������ "�T6^6F�X�j�a��r�ϔ�����	��������t����>0 ����y��
SM #\'�	��X��	��r!��h�z�@��Ugy�3�� ������"4�FX�����A�Z��nn���		������ //&/8/J/\/n/�/ �/�/�/�/�/�/�/?"?2<�2?V?h?z?�? �?�?�?�?�?�?
OC �~(O����O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_@?oo,o>oPo boto�o�o�o�oOJO <O`OrO:L^p ������� � �$�6�H�Z�l�~��� �_��Ə؏���� � 2�D�V�h�z��o���� 0��
��.�@� R�d�v���������Я �����*�<�N��� r���������̿޿� ��&�8ϴ���P�ʟ ܟ���������� "�4�F�X�j�|ߎߠ� �����������h�0� B�T�f�x������ ����@�r�d�-��Ϛ� b�t������������� ��(:L^p �������  $6HZl~� �����4�F�X� / 2/D/V/h/z/�/�/�/ �/�/�/�/
??.?@? R?d?v?��?�?�?�? �?�?OO*O<ONO`O ��xO�//�O�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4o�?Xojo|o�o�o �o�o�o�o�ohO�O �OU�O�O���� �����,�>�P� b�t���������Ώ�� <o��(�:�L�^�p� ��������ʟ&�� \n�H�Z�l�~��� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
��.�@� R�d�vψ������� ,�>���*�<�N�`� r߄ߖߨߺ������� ��&�8�J�\︿�� ������������� "�4����ϴ�}����� ����������0 BTfx���� ���d�>P bt������ �N�/
/������p/ �/�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�? �?�?�?"�?�?O O 2ODOVOhOzO�O�O�O ,//�OB/T/f/._@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�?�o�o�o�o�o &8J\�O�O �O� __���� "�4�F�X�j�|����� ��ď֏�����0� �oB�f�x��������� ҟ�����v?�2� ���������ί� ���(�:�L�^�p� ��������ʿܿ�J� �$�6�H�Z�l�~ϐ� �ϴ�����T�F���j� |���V�h�zߌߞ߰� ��������
��.�@� R�d�v������� ������*�<�N�`� r���������(�:� &8J\n� ������� "4FX��j�� �����//0/ B/��g/Z/�������/ �/�/�/??,?>?P? b?t?�?�?�?�?�?�? �?OOr:OLO^OpO �O�O�O�O�O�O�O _ |/n/_�/�/�/~_�_ �_�_�_�_�_�_o o 2oDoVohozo�o�o�o �o�o0O�o
.@ Rdv���_:_ ,_�P_b_*�<�N�`� r���������̏ޏ�� ��&�8�J�\�n��� �o����ȟڟ���� "�4�F�X�j������ �� ������0� B�T�f�x��������� ҿ�����,�>Ϛ� b�tφϘϪϼ����� ����(ߤ���@ߺ� ̯ޯ�߸������� � �$�6�H�Z�l�~�� �����������X� � 2�D�V�h�z������� ����0�b�T�xߊ� Rdv����� ��*<N` r������� //&/8/J/\/n/�/ �/���/�/$6H? "?4?F?X?j?|?�?�? �?�?�?�?�?OO0O BOTOfO��O�O�O�O �O�O�O__,_>_P_ �/�/h_�/�/?�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $�OHZl~� ������X_�_ |_E��_�_z������� ԏ���
��.�@� R�d�v���������П ,���*�<�N�`� r����������߯ү L�^�p�8�J�\�n��� ������ȿڿ���� "�4�F�X�j�|ώ�� ������������0� B�T�f�x���毐�
� �.�����,�>�P� b�t��������� ����(�:�L���p� ��������������  $�߲ߤ�m���� ������  2DVhz��� ����T�
/./@/ R/d/v/�/�/�/�/�/ �/>?�/t��`? r?�?�?�?�?�?�?�? OO&O8OJO\OnO�O �O�O�O/�O�O�O_ "_4_F_X_j_|_�_�_ ??�_2?D?V?o0o BoTofoxo�o�o�o�o �o�o�o,>P bt�O����� ���(�:�L��_�_ �_���_oʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � |2�V�h�z������� ¯ԯ���
�f�/�"� ��������������п �����*�<�N�`� rτϖϨϺ�����:� ��&�8�J�\�n߀� �ߤ߶���D�6���Z� l�~�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt����߽�*� �(:L^p ������� / /$/6/H/��Z/~/�/ �/�/�/�/�/�/? ? 2?�W?J?����? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O�O �O�O_b/*_<_N_`_ r_�_�_�_�_�_�_�_ l?^?o�?�?�?no�o �o�o�o�o�o�o�o "4FXj|�� �� _����0� B�T�f�x������_*o o�@oRo�,�>�P� b�t���������Ο�� ���(�:�L�^�p� �������ʯܯ� � �$�6�H�Z����r� ����ؿ���� � 2�D�V�h�zόϞϰ� ��������
��.ߊ� R�d�v߈ߚ߬߾��� �������0謹 ��ο���������� ��&�8�J�\�n��� ������������H� "4FXj|�� �� �R�D�h�z� BTfx���� ���//,/>/P/ b/t/�/�/���/�/�/ �/??(?:?L?^?p? �?��?�?&8 O O$O6OHOZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_�/z_�_�_�_ �_�_�_�_
oo.o@o �?�?Xo�?�?�?�o�o �o�o*<N` r������� ��p_8�J�\�n��� ������ȏڏ�Hozo lo5��o�oj�|����� ��ğ֟�����0� B�T�f�x��������� �ү����,�>�P� b�t��������Ͽ¿ <�N�`�(�:�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~�گ �ߴ���������� � 2�D�V�h��ֿ���� ������
��.�@� R�d�v����������� ����*<��` r������� p���]���� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/D�/?0? B?T?f?x?�?�?�?�? �?.�?�?dv�PO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_?�_�_�_ o o$o6oHoZolo~o�o O�?�o"O4OFO  2DVhz��� ����
��.�@� R�d��_��������Џ ����*�<��o�o �o���o�o��̟ޟ� ��&�8�J�\�n��� ������ȯگ���� l�"�F�X�j�|����� ��Ŀֿ���V��� ������xϊϜϮ��� ��������,�>�P� b�t߆ߘߪ߼���*� ����(�:�L�^�p� �����4�&���J� \�n�6�H�Z�l�~��� ������������  2DVhz��߰ ����
.@ Rd�������� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?�J?n?�? �?�?�?�?�?�?�?O "O~GO:O����O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_R?o,o>oPo boto�o�o�o�o�o�o \ONO�orO�O�O^p ������� � �$�6�H�Z�l�~��� ����o؏���� � 2�D�V�h�z����o ՟0B
��.�@� R�d�v���������Я �����*�<�N�`� ��r�������̿޿� ��&�8�JϦ�o�b� ܟ� ���������� "�4�F�X�j�|ߎߠ� ������������z� B�T�f�x������ ���������v� ��� �Ͼφ����������� ��(:L^p ������8�  $6HZl~� ���B�4��X�j� 2/D/V/h/z/�/�/�/ �/�/�/�/
??.?@? R?d?v?�?��?�?�? �?�?OO*O<ONO`O rO��O�O//(/�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4oFo�?jo|o�o�o �o�o�o�o�o0 �O�OH�O�O�O�� �����,�>�P� b�t���������Ώ�� ��`o(�:�L�^�p� ��������ʟܟ8j \%���Z�l�~��� ����Ưد���� � 2�D�V�h�z������� �¿���
��.�@� R�d�vψϚ����ϲ� ,�>�P��*�<�N�`� r߄ߖߨߺ������� ��&�8�J�\�n�ʿ ������������� "�4�F�X�����p��� ���������0 BTfx���� ���,��P bt������ �/`�����M/���� �/�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�? �?�?�?�?4�?O O 2ODOVOhOzO�O�O�O �O/�O�OT/f/x/@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�?�o�o�o�o &8J\n� �O�O�_$_6_�� "�4�F�X�j�|����� ��ď֏�����0� B�T��ox��������� ҟ�����,��� �u�������ί� ���(�:�L�^�p� ��������ʿܿ� � \��6�H�Z�l�~ϐ� �ϴ�������F��� |�����h�zߌߞ߰� ��������
��.�@� R�d�v������ ������*�<�N�`� r�������$����:� L�^�&8J\n� ������� "4FXj|�� �����//0/ B/T/�������/��
 �/�/�/??,?>?P? b?t?�?�?�?�?�?�? �?OO(O�:O^OpO �O�O�O�O�O�O�O _ _n/7_*_�/�/�/�_ �_�_�_�_�_�_o o 2oDoVohozo�o�o�o �o�o�oBO
.@ Rdv����� L_>_�b_t_�_N�`� r���������̏ޏ�� ��&�8�J�\�n��� ���� ȟڟ���� "�4�F�X�j�|��
� �ů �2�����0� B�T�f�x��������� ҿ�����,�>�P� ��bφϘϪϼ����� ����(�:ߖ�_�R� ̯ޯ�������� � �$�6�H�Z�l�~�� ������������j� 2�D�V�h�z������� ��������t�f��� �߮�v����� ��*<N` r�����(�� //&/8/J/\/n/�/ �/�/ 2$�/HZ "?4?F?X?j?|?�?�? �?�?�?�?�?OO0O BOTOfOxO��O�O�O �O�O�O__,_>_P_�b_�%�$SBR2� 1�%�P �T0 � �	C�/�' �_�_�_�_ oo&o8oJo\ono�o�o�o�o�Q�o�_�o '9K]o� ������o��o #�5�G�Y�k�}����� ��ŏ׏�����1� �U�g�y��������� ӟ���	��-�?�"� c�F���������ϯ� ���)�;�M�_�q� T���x���˿ݿ�� �%�7�I�[�m�ϑ��φ�~i_������� �'�9�K�]�o߁ߓ� �߷����ظ���
�� .�@�R�d�v���� ������������*�<� N�`�r����������� ����&
��\ n������� �"4FX<f �������/ /0/B/T/f/x/�/n �/�/�/�/�/??,? >?P?b?t?�?�?�?�? �/�?�?OO(O:OLO ^OpO�O�O�O�O�O�O �O�?_$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ o o_DoVohozo�o �o�o�o�o�o�o
 .@R6ov��� ������*�<� N�`�r���h����̏ ޏ����&�8�J�\� n�����������ڟ� ���"�4�F�X�j�|� ������į֯��̟� �0�B�T�f�x����� ����ҿ������ >�P�b�tφϘϪϼ� ��������(�:�� ^�p߂ߔߦ߸����� �� ��$�6�H�Z�l� Pߐ����������� � �2�D�V�h�z��� ������������
 .@Rdv��� �����*< N`r����� ��/�&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?4?/X?j?|? �?�?�?�?�?�?�?O O0OBOTO8?J?�O�O �O�O�O�O�O__,_ >_P_b_t_�_jO|O�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�_�o �o $6HZl ~�������o � �2�D�V�h�z��� ����ԏ���
��  �@�R�d�v������� ��П�����*�<� N�2�r���������̯ ޯ���&�8�J�\� n���d�����ȿڿ� ���"�4�F�X�j�|� �Ϡϲϖ�������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� �����������:�L� ^�p������������� �� $6�,�l ~�������  2DVhLv ������
// ./@/R/d/v/�/�/~ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �/�?OO&O8OJO\O nO�O�O�O�O�O�O�O �O�?"_4_F_X_j_|_ �_�_�_�_�_�_�_o o0o_Tofoxo�o�o �o�o�o�o�o, >PbFo���� �����(�:�L� ^�p�����x��ʏ܏ � ��$�6�H�Z�l� ~�������������� � �2�D�V�h�z��� ����¯ԯ�ʟܟ� .�@�R�d�v������� ��п�������&� N�`�rτϖϨϺ��� ������&�8�J�.� n߀ߒߤ߶������� ���"�4�F�X�j�|� `ߠ����������� �0�B�T�f�x����� ����������, >Pbt���� ����(:L ^p������ � //�6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?D?(/h?z?�? �?�?�?�?�?�?
OO .O@OROdOH?Z?�O�O �O�O�O�O__*_<_ N_`_r_�_�_zO�O�_ �_�_oo&o8oJo\o no�o�o�o�o�o�_�o �o"4FXj| ��������o �0�B�T�f�x����� ����ҏ�����,� �P�b�t��������� Ο�����(�:�L� ^�B���������ʯܯ � ��$�6�H�Z�l� ~���t���ƿؿ��� � �2�D�V�h�zό� �ϰ��Ϧ�����
�� .�@�R�d�v߈ߚ߬� �����������*�<� N�`�r������� ��������
�J�\� n��������������� ��"4F*�<�| ������� 0BTfx\� �����//,/ >/P/b/t/�/�/�/� �/�/�/??(?:?L? ^?p?�?�?�?�?�?�? �/ OO$O6OHOZOlO ~O�O�O�O�O�O�O�O _�?2_D_V_h_z_�_ �_�_�_�_�_�_
oo .o@o$_dovo�o�o�o �o�o�o�o*< N`rVo���� ����&�8�J�\� n��������ȏڏ� ���"�4�F�X�j�|� ������ğ������� �0�B�T�f�x����� ����ү���ڟ�,� >�P�b�t��������� ο����(��6� ^�pςϔϦϸ����� �� ��$�6�H�Z�>� ~ߐߢߴ��������� � �2�D�V�h�z�� p߰���������
�� .�@�R�d�v������� ��������*< N`r����� ����&8J\ n������� �/"/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?8/x?�?�? �?�?�?�?�?OO,O >OPObOtOX?j?�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�O�O�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�_�o  2DVhz� ������
��o .�@�R�d�v������� ��Џ����*�<� N�