��   D�A��*SYST�EM*��V9.1�0170 9/�18/2019 A 
  ����CELLSE�T_T  � w$GI_ST�YSEL_P �7T  
7ISO:iRibDiTRA�R|��I_INI; �����bU9A�RTaRSRPNSS1Q23U4567y8Q
TROBQ?ACKSNO� �)�7�E� S�a�o�z�2 3 4 5* 6 7 8aw.n&GINm'D�&� �)%��)4%��)P%���)l%SN�{(O�U��!7� OPT�NA�73�73.:BP<;}a6.:C<;CK;�CaI_DECS�NA�3R�3�TR�Y1��4��4�PTHCN�8D�D>�INCYC@HG��KD�TASKOK�{D�{D�7:�E �U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbH<aRBGSOLA�6�VbG�S�MAx��Vp��Tb@SEGq��T��T�@REQ �d�drG�:Mf�G�JO_HFAUL��Xd�dvgALE@� �g�c�g�cvgE� x�H�dvgNDBR�H<�dgRGAB�Xt�b���CLMLI�y@   �$TYPESIN�DEXS�$$C�LASS  ����lq�����apVERSION�ix  ��Z�$'61�r���p��q�t+ �UP0 �x�Style Se�lect 	  ���r�uReq. _/Echo���y�Ack�s�sI?nitiat�p�r��s�t@�O�a�dp���	��  ��U��������:q�������q��s�Option b�it A��p�B�����C�Deci�s�cod;��zTryout mL���Path se}gJ�ntin.��II�yc:��Ta�sk OK��!�M�anual op�t.r�pAԖB�ޟԖC�� dec�sn ِ�Rob�ot inter�lo�"�>� isSol3��C��i/�<"�z�ment���z�ِ����_�sta�tus�	MH ?Fault:��ߧOAler�#����p@r 1�z �L��W�i�{��$�; LE_COMN�T ?�y�   ��䆳�Ŀֿ� ����0�B�T�g�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼�������������U��9r��   ���ENAB  ���u�����x���ꐵMENU>���y��NAME ?=%��(%$*4��� D��p2�k�V���z��� ����������1 U@Rdv��� ����*< u`������ ��/;/&/_/J/f/ n/�/�/�/�/�/?�/ %??"?4?F?X?j?�? �?�?�?�?�?�?�=