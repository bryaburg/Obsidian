��   ?3�A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����MN_MCR�_TABLE �  � $MA�CRO_NAME� %$PRO�G@EPT_IN�DEX  $OPEN_IDa�ASSIGN_T�YPD  qk$MON_NO}�PREV_SUB�y a $USER�_WORK���_�L� MS�*RT�N  _&S�OP_T  �� $�EMG�O��RESE�T�MOT|�H�OLl��12��STAR PD�I8G IAGBzGC�TPDS��REL�&U�s �� �EST�x��SFSP�C���C�C�NB��S)*$8�*$3%)4%)5%)6�%)7%)S�PNS�TRz�"D�  ��$$CLr   O����!������ VERSIO�N�(  ��Z�:LDU�IMT  ���� ����$MAX�DRI� ��5
��$.1 �%� � d%�Open Gri?pper 2����%  RIPP� pfZ?���"  �!���q0Clos�eQ?d?v4CLOS�E�?�?�0�4Re�lax hand3 1�?�6 )OOO�9�#q0M2B�?@1O�OUO�4 qD�3 ~O�O__�8�GH �O�Oo__�3oFh_ �_d_�_�[�3�5�_o �_=o�_�_so"o�oFo Xo�o�o�o�o�o9 �oIo0�T� x����5��� k����>�P���׏ ������1���U��� P���L���p������� �ʟܟ�c����6� H���l�ͯ󯢯��)� دM������2����� h�z�￞��¿Կ!� [�F��.�@ϵ�d��� �Ϛ���!���E���� {�*ߟ�N�`ߚ��ߖ� ����A���Q�w�&� 8��\��������pp3-�?�����+� x�'���K�]������� ����>��b# �G��}�� (��^p[�C U�y���$/6/ �Z/	//�/?/�/c/ u/�/�/�/ ?�/�/V? ?z?�?;?M?�?q?�? �?�?O�?@OROOO �O7O�O[OmO�O�O�O _�O�ON_�Or_!_3_ �_�_i_�_�_�_o�_ 8o�_�_3o�o/o�oSo eo�o�o�o�o�oF �oj+�O�� ����0���f� x�c���K�]�ҏ���� ����,�>��b��#� ��G���k�}������ (�ן�^������C� U�ʯy����$�ӯ H�Z�	����?���c� u����� �Ͽ�V� �z�)�;ϰ���q��� �ϧ����@����;� ��7߬�[�m��ߑ�� �����N���r�!�3� ��W���������� 8�����n���k���S� e�����������4F ��j+�O�s ���0��f ��K]��� ��,/�P/b//#/ �/G/�/k/}/�/?�/ (?�/�/^??�?1?C? �?�?y?�?�?�?$O�? HO�?	OCO�O?O�OcO uO�O�O_ _�O�OV_ _z_)_;_�___�_�_ �_�_o�_@o�_ovo �oso�o[omo�o�o �o�o<N�or!3 �W�{���� 8���n������S� e�ڏ��������4�� X�j��+���O�ğs� �������0�ߟ�f� ���9�K���ү���� ����,�ۯP����K� ��G���k�}�򿡿� (�׿�^�ς�1�C� ��g����ϝϯ�$��� H���	�~ߐ�{ߴ�c� u��ߙ�����D�V� �z�)�;��_���� �������@����v� %�����[�m����� ����<��`r!3 �W�{�� 8��n�AS ������4/� X///S/�/O/�/s/ �/�/�/?0?�/�/f? ?�?9?K?�?o?�?�? �?�?,O�?PO�?O�O �O�O�OkO}O�O�O_ �O�OL_^__�_1_C_ �_g_�_�_�_�_$o�_ Ho�_	o~o-o�o�oco�uo�o�o�dOVE��o�oN.r?x �ETI+=� pV�AL�� $CUp��� pR_A�@�  $��z��qR��   a	W�i�ޏ�� Ϗ� ACH��͏B�� pD fk�   !	�o0�������П� TR*��	��rL.�3��pER���n�F p_V���O�K��]�ү)�ROï�� � ����5��� $<'�`� _DA�%���� pCMD��Ŀ a������S�AT��(���^��dUR_�SόϬ���P����sJ�����cq�ϵ�*ߍ�R��T߷�ߊ��e@�߸��oy��$MA�CRO_MAXN�U  �d��� p���SO�PENBL ��������o��A��b�PDIMS�K����Y�S�Uc�u�TPDSB�EXR�_tq�U� ���n����