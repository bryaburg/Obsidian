��   v��A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@ � &�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	>4SUSRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  ��Z�$'2 ��\���R	 /,��?���aa1`jbed`a�����[`�� �`dc�o��
 ��a�o�o�o%7 �o\n�� ��E����"� 4��X�j�|��������ď�)/SOFT�P�@/GEN�1?�current=�menupage,1422,1ŏ �%�7�ƏT�m���� ����ǟV�����!� 3�E�ԟi�{������� ïR�d�����/�A� S��w���������ѿ��� TPTX��l����a`� s縄�$/�softpart�/genlink�?help=/m�d/tp�.dg ޿xϊϜϮ�g����� ����,߻�P�b�t� �ߘߪ�9߻������ �(�:���^�p���X������a�fq�b�b�� ($R������6�!�Z��i  ada��c�������N��k
��adJ��aJ�  �8J�PJ������4`�~�~��b���`�  ���H GpO��K#J��FF��I�:c�B 1�)hR \���_�� ;REG VED?����wholem�od.htm�	s�ingl�do�ubtri�pbrows3b�i{�W �����"/��|��dev.s��lo/� 1r,	t �/A�//K/�/�/?��/5?G?Y?k?}?�?� `�?�?�?�?O O*O<ONO`OjF2P�? �O�OqO�O�O�O�E�	 �?�?_/_A_S_e_w_ �_�_�_�_�_�_�_o o+o=oOoao/'yoso �o�o�o�o�o�o 1CUgy��� ����? �2�D�V� h�z��������O� ��Ǐُ.�@��O	_� ��������П˟ݟ� ��%�7�`�[�m�� �������oկϯ��� !�3�E�W�i�{����� ��ÿտ�����/� A��|ώϠϲ����� �������B�T�#� 5ߊߜ�S�e�K����� ���,�'�9�K�t�o� ������������ �߯1�+�Y�k�}��� ������������ 1CUgy��k� ��� 2DV hzuߞ��� ����ߧ@/;/M/_/ �/�/�/�/�/�/�/�/ ??%?7?`?[?m?;� �?�?�?�?�?�?�?O !O3OEOWOiO{O�O�O �O�O�O�O�O�4_F_ X_j_|_�_�_�_�_�_ ��_o�_�_BoTobj��$UI_TOP�MENU 1�-`�aR �
d�aQ)*default_� ]*leve�l0 *[	 �o�0�o�o�o	r�tpio[23]��8tpst[1�=xY�o�o�=�h58e01_l�.png��6m�enu5�y�p�q1!3�z�r�z�t4�{��q��?�f�x����� ����RT�������1�C�҄prim�=�qpage,1422,1J����� ����˟֏���%��7�I�ؖ^�class,5R�������h��ϯڔf�13֯@��0�B�T�ۓ^�53p�������ƿؿ
ۓ^�8��%�7� I�[�ڟϑϣϵ�����Y�`�a�o��m�Ιq�;�mCvtyxN}6Hqmf[0P�N�	��c[164=w��59=x�q)�[�&�tc8�|�r2��} Q����w�{��O�� ����� ��$�o�H��Z�l�~�����Q�c�80������	-`�r�22gy��� >p���	-� ���n����e�w�1���//*/</�7�^�ainedi	�s/�/�/�/�/2��config=single&^�wintpj��/? ?*?<?����r?!ٙ�gl[55�ٕSߐ�?�;Ip�08�ݔ07A6=y�?�5���62,O[I�?	OoO�z��z�4s�x�O�� �x� �B�Q�*_<_N_ `_r_�_3��_�_�_�_ �_o�_&o8oJo\ono�o�o�!;�$dou�b�%oc�13~�&odual�i38��C,4�o�o�o9�o �n�o�ax��#o��������%3B.=_!g�Q�b8"� z�������\ԏ����
���+:6��i48,2Q��b]������ ]?ҟ�/�UE������s���_����G�u��:���"�f7 .�ݣB�Or��J�\�6G�u7������ÿտ翮��27 ��)�;�M�_�q� �ĀU�����������!�1�/�A�S�e�w� ��߭߿������߄� �+�=�O�a�s��� �������������6
�?�Q�c�u����$��74�����������C���6�	TPTX[209�<aAY2+H,���BY1�8t?Ht���a
t0�2��aA��=�DtvB��O�L_��0��Li�S=�treeview�#�X�3��`�381,26�o//A/S/�w/ �/�/�/�/�/`/�/? ?+?=?O?�o�
��o`%���?�?�?�Ar?">1`��?"2��GO YOd?v?�_�.E-��O �O�OxO��@�O0OC_U_g_��6�OF�'_n_ �_�_�_8�_���_�S �_Qocouo$vo�o� �o#�oS�o�o 1CUz�os�� ����
��y�3� Z�l�~��������/؏ ���� �2���V�h� z�������?���� 
��.�@�ϟd�v��� ������M������ *�<�˯N�r������� ��̿[����&�8� J�ٿnπϒϤ϶��� wo�o�ϭo"߉'�E� W�i�{ߎߟ߱���1� ������/�A�S�e� w�9������������ �e�>�P�b�t����� '����������� :L^p���5 ��� $�H Zl~��1�� ��/ /2/�V/h/ z/�/�/�/?/�/�/�/ 
??.?����d?߈? �ߍ�?�?�?�?�?O O)O�?5O_OqO�O�O �O�O�O�O��_&_8_ J_\_n_�_�/�_�_�_ �_�_�_�_"o4oFoXo jo|oo�o�o�o�o�o �o�o0BTfx ������� �,�>�P�b�t����� '���Ώ������� :�L�^�p�����C?U? ʟy?�UO�O�#�5� G�Y�k�~�������ů ׯ�����1�C�_ z�������¿Կ�� 
��.�@�R�d��� �ϬϾ�����q��� *�<�N�`���rߖߨ� ����������&�8� J�\�n��ߒ����� ����{���"�4�F�X� j�|�������������������*def�ault؞*?level8a����Y�w�! t?pst[1]�	��y�tpio[#23���u�d��,>menu7_l.pngAM^13cp5xh]�[4�u6c p���	//-/?/�� c/u/�/�/�/�/L/�/��/??)?;?M?�"�prim=^page,74,1R?@�?�?�?�?�?�"f6�class,13 �?OO0OBOTO�?�25ZO�O�O�O�O�O�#�<~O_$_6_H_Z_]?o218v?�_�_�_�_�_�O�26�_o-o�?oQocoB�$UI�_USERVIE�W 1�����R 
�A�jo䒞o�o=m�o �o	-?�ocu ���N���� ��o$�6�H������ ����ˏn����%� 7�I��m�������� `�ԟ�X�!�3�E� W�i��������ïկ�x�����/�A���*zoomT�ZOOMIN�S�� ��̿޿�ϥ�&�8� J�\�n�ϒϤ϶������<*maxre�sn�MAXRES ���ω�R�d�v߈ߚ� =߾���������*� <�N�`�r�߃��� �������&�8��� \�n�������G����� ������3A�� |����g�� 0B�fx� ��Y���Q/ ,/>/P/b//�/�/�/ �/�/q/�/??(?:? �K?Y?k?�/�?�?�? �?�? O�?$O6OHOZO lOO�O�O�O�O�O�? �O�O	_{OD_V_h_z_ �_/_�_�_�_�_�_
o �_.o@oRodovoa