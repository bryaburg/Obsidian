��   8��A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����DCSS_I�OC_T   �P $OPER�ATION  $L_TYPB7IDXBR1H[ �S2]2R �$�$CLASS  �������Pz��P� VERS?��  ��Z�$' 2 ��P @+ ������ $B �
��� ���"����A����:G��F�����:@����b��T ���38��b  	$
/ �&!�J�B/�������2 ������ O(�!&!!��R%�! &!�:%R%�!�%�%� :�!5A?S?e?w?�? �?�?�?�?�?�?OO +O=OOOaOsO�O�O�O �O�O�O�O__'_9_ K_]_o_�_�_�_�_�_ �_�_�_o#o5oGoYo ko}o�o�o�o�o�o�o �o1CUgy��������_C_CCL ?���  	All param���
Base��Pos./Sp�eed chec�k(�Safe I�/O connect�}R��� �X2�D�V�SIi�@{� �����!�3�J�W� i�{�������ßڟ� ���"�/�A�S�j�w� ��������ѯ���� �+�B�O�a�s����� ����ҿ߿���'� 9�K�b�oρϓϪϷ� ���������#�:�G� Y�k߂ߏߡ߳����� ������1�C�Z�g�y�������ކO �����%�N�I�[�m��������at pi���������� =8J\���� ����"4 ]Xj|���� ���/5/0/B/T/ }/x/�/�/�/�/�/�/ ???,?U?P?b?t? �?�?�?�?�?�?�?O -O(O:OLOuOpO�O�O@�O�O�O�O_��N�  {��	_��;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{� ���������SIh���Ob����� ����ӏΏ����� (�:�c�^�p������� ��ʟ�� ��;�6� H�Z���~�����˯Ư د��� �2�[�V� h�z�������¿�� ��
�3�.�@�R�{�v� �Ϛ��Ͼ������� �*�S�N�`�rߛߖ� �ߺ��������+�&��1�P%_�W�SF'DI10�y�2�y�I3��y�4��y�5��y�6��y�7��y�8 �G�3�E�W�n�{��� ������������ /FSew��� ����+= Ofs����� ��//'/>/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?^?k?}? �?�?�?�?�?�?�?O O6OCOUOgO~O�O�O �O�O�O�O�O__-_ ?_V_c_u_�_�_�_�_ �_�_�_oo.o;oMo _ovo�o�o�o�o�o�o �o%7N[m ������� �&�3�E�W�n�{��� ����ÏՏ����� /�F�S�e�w������� ��֟�����+�=�$H�Z�Od�v�O~ ���� ����&�`�Q�c� ��������ԿϿ�� ��)�;�d�_�qσ� �ϧϹ��������� <�7�I�[߄�ߑߣ� ����������!�3� \�W�i�{������ �������4�/�A�S� |�w������������� +TOas ������� ,'9Kto�� ����/�/#/ L/G/Y/k/�/�/�/�/ �/�/�/�/$??1?C? l?g?y?�?�?�?�?�? �?�?	OODO?OQOcO �O�O�O�O�O�O�O�O __)_;_d___q_�_ �_�_�_�_�_�_oo�<o7oIo[o�ox�SIz����VOFFno�FENCE�oEXEMG�o�o�c�NTED�OP�oqAUTOT��[s���a�MCC|pCS�BP�
POSSPD_ENB�j�CONF_OK��~F_IPAR_�CR�z�g����~��o�q_�o;��o�`�'�DIS�|C_�r_`��y 