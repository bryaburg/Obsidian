��   �A��*SYST�EM*��V9.1�0170 9/�18/2019 A 	  ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTT  &F/�� $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STSTOP�_TPCHG �V LOG_P NT��N�  6 C�OUNT_DOW�N�$ENB_�PCMPWD� �$DV_� IN�� $C� CR5E��A RM9� =T9DIAG9(|�LVCHK >FULLM/��YXT�CNTD��MENU�A�UTO+�FG_wDSP�RLS��U�BURYBAqN�!eENC/�  CR�YPTE ����$$CL(  ? ���K!��� T @ V� ION�H(; �Z��$DCS_COMD?���O%�H e^z'_� �-W�(WS  J*�� L ��&�A91�"K!�	 
 $R!��=?$?2?H? V?l?z?�?�?�?�?�? �?�?
O O.ODO<#'WSUP� �*�FOXO�#FxO�O�O>��  �L�A���_ � �� �V�[t&��j
���D�O`_��W�_��;!�U�_cGLU�GH 1K) ; �)�_�_ 	oo-o?oQocouo�o �o�o�o�'�_�o�o !3EWi{�� ���o����/� A�S�e�w��������� ������+�=�O� a�s���������͟܏ ���'�9�K�]�o� ��������ɯ؟د�� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� �������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q����������� ��%�7�I�[�m�� �������������� !3EWi{�� �����%