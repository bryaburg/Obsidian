��   6�A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	  /GR�P:� $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2� RING,��<$]_d��REL3� 1  	��CLo�: � �A�X{  $PS_��TI���TI�ME �J� _gCMD��"FB��VA �&CL_OV��� FRMZ�$DmEDX�$NA� �%�CURL��W���TC�K�%�FMSV��M_LIF 	��'83:c$�-9_09:_��=�%3�d6W� �"�PCC�OM��FB� M��0�MAL_�E�CI�P:!o"DTYkR_|"�5:#N�1END�4��^o1 l5M����PL� W� ��STA:#T�RQ_M��� K$NiFS� uHYsJ� �hGI�JI�JI�D���$�ASS> �����A����>�@VERSI� �G�  �wZ�$S 1�H� ����N ��>_)_b_MV���" ���X��mJ ?<���:��(_ �_t_�_H]P�X	oPU��A$om
� ��q m�m���#���X�e��oroo7l�o�o��o�o�`����5��  (�g�� uggB@v 'w�oooXC|���do�����=gL����?����@��D�V�h�z� ������ԏ���
�] �E5�C�-�c��D  2������� ʟܟ� ��$�6���<��`�r����������̯ޯ���&�a|( mZ�i~�i�����ƿ ��ÿ��� ��D�/ϰh�S�xϞ��$4 �1\��H��G�0�H��oN���K���Hx�}�O�!��POΔO���F��H?𧻓K���ʯFC� "ߤ|���畒�ƥE���Gb@���u�½S�����zQ�mP�:QCF�ƠI��K�~�}��A����|�H���G�9�H�}���"H}l��T� ܉����\��o��L�7��Tȿ2DT�Cw:����  c�����n �W�T��W:������.�ta�>A�UY����7j.�������b1�X�,>7A��V5ߡ��3�.�>I� ��s��Aj��f>�Qx@���P�^Q�~ ����%�@�1LOSEQ����������� Hг�	�}�Ń��O���S
��Bp�}:޳�p����u����<��O�d�Bp�?�.�@�_A�9ۉ��v4>����B~����5;��"��PLACE� e I�C�LL�LEF�T!��R�Ǩm���C
�A#���un.�k(�A�U:��B��Al�����g9(�or�A���.�����pA�|���YȽ��"�A��@� ��������X���K�r��A���A�^Xb���f����B�a�.�B��A��F��W�ɿ������RB���f�h_B�x���A���>�A�3_A�ێ�"����RIGH���(�d���r�@'B8����@�@���]���B����)�B7����|@�F��^�B�Q�o��C>�}rA�5�?Ɛ@!�������N��"�GRIPP��0OPE�@5/(���`�r2t�B�s����$@�}���6CB��c��B2l�B�sw`��8@W}��v �z �.����2@A��@��>������v��(��/ $gy+��R�ʫ �F�WN��R��V�^Z�[^�a>ۅ�J���T��O�B@�7��S^��0���p�@][�?<3��?[+�A�A�o?4�x�/�"/�?/F/6�FӒ������D�@���������T�>?����	�����@��,<�½�V.������BAM��>����@99=1(��?�4���1����琠��mX���+@�2��ؓ�0��?��:�ێ��� ��@�Kߘ½Uqf>��z��;3AF��%>��A@z��=&��NO�1�ufOxO�O�0�I��^-A�7����a@�W����LB�f_��n�A�����-@��A�uwB�q��;�=�@�Y����@��i�?��A�
//�?�?R[�Qbr�Z��������������oB�5��o|���GH��uĿ��.�/�B�ˑ7�?���A����������,�A��@8�6�_`�/D_h���	K��X�����.�N��_B`2���W��������d���BY�&N�4]���q�A�.+X>���@�&~>a�\�o`�d�_xo]PT����\���]���B>A'��U�E���|��\*���l���>'���V2 ���s{sa7���&��A���>�l��@/�= �&N �2�D�V��	���������X�>A	���Uu[��Q���������c��>-O��V��z��4�&N2���?D@�@�2�;>�OhA/�?�4��_�1�C���S:�����Bu_�.����Ң�9��C4V�.������B �4�-�<ɻ�@ �:�!C4T!������?�7@���8>��a@��>J�g|����T�3������4����P�
��{�p�Bv��o��տ��p���+C�|*�Bt'.�1�OO����AU��>Q(N@�?IL><Ύ�`貟ğ֘��������������ن�{iWB��/>o���������@��p�|�B��P�^ e��a���A2�>��@��f>��]�o���Ӛ��F���|�Ñ������@p�{��.¾�h�O����ۮ����@ņ�|X��¾�������n�gA90�>�<x@����A�8ܜ?.�@�қ˽�b��r�������z��;[�>-f��V�x���&�+�Q�
��C1�A)�>�o�A��<�^�ο�����V�U�F����P��{�@��i�d7���^W~�a�rE�5��֡@^�����S��f>���@$e��?��w?[O3Au�"�����޿�����;�2�UОߤЌ��$P�LCL_GRP �1�@����?� D�sa��  ��x�O?r����:���8� J�5�n�Y��}���������� 