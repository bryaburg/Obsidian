��   �=�A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����EIP_CF�G_T   �� $VENDO�R  $DE�VTYPE>PR�DCODIREV�ISION>FA�ST_UDP �5 KEEP_IO�_AnSCNpO�PT` Sp $L�OADED� �C�C� IG�ED_wMOD�NET��EXPLCIT_�MS�$HIG�H_SPEE�$EN8021p�DSCP� Hp ��� SPARE�� &ONN.� | $HOS�� !B SC9E�NABL$S�TATN _SZ��S^TOAPI�OTrIgA��R]V�BW&MjoD&SC.�  7�C`XQ�[XX_���X_��[ kqRs)%'FLA�7MUL�TR�� gC_O�["TOD&�ICi �AS��Z 'EC{#�#TI�MVCN� Z�&P�AT  @$�IDA_FORM�A��!�&� �"9"F�IG^�"2�+�!��$ANALOG�I�   4O�U� 8FM�$�Q�(O8�$$C�LASS  ����e1��.��.�Z0VER_c7�  �Z��$'0 �8. d*���� ���0��?��0���7/ ���4( 2�;@� p!
11.2�00.1.1�����+ �=Oas � �!ConnectionB(CO�5�1_D gD�:�!�3   h;{{Yx�A@�  � �\ !��P�0p3I2HO��bENMzE�O��3I3_1_C_�Og_
_<@4q_�_�_V_�_z_<@5�_o#o�_Go�_<@6Qo�o�o6o�oZo<@7�o�o�o'�o<@81as�:<@9������<@A�A�S��w��<@B����Ïf����<@C�!�3�֏W���<@Da�����F�ǟj�<@Eџ����7�ڟ<@FA�q���&���J�<@G���󯖯���<@H!�Q�c����*�<@I����ӿv�����<@J�1�C��g�
�<@Kqϡϳ�V���z�<@L���#���G���<@MQ߁ߓ�6߷� Z�<@0���ߖߨ�)���nO1�a�s���:�<@P����������<@Q�A�S���w��<@R������f��� ��<@a0#����Y��nTa��F�j<@U��7�<@VAq�&�J<@W����/
�5A3_K/]/ / �/$/6!�_�/�/p/�/ �/6!�_+?=?�/a?? 6!oo�?�?P?�?t?6! �oOO�?AO�?�1O {O�O0O�OTO�1��O`�O�O!_�O�0401_@\_n__�_5_GP1�_@�_�_�_o�_GP2o <oNo�_rooGP:/�o �o`o�o�oFQ�/- �oQ�oFQ?��@ �dFQ�?���1� �FQ�?k�}� ���D� FQjOۏ폐����FQ��OK�]� ���$��05 J_��͟p�񟔟���_ +�=���a����*o�� ��P�ѯt����o�� ��A�䯦�
{���0� ��T���z�����!� Ŀ���[�m�ϑ�4� ��Z����π�ߤϦ� ʏ;�M���q�ߦ�:�@�߽�`��߄��06�� �-���Q������� ��@���d�ኯ��� ��1������k�}� ����D��j���������$EIP_SC �2����. @����� K�������A@]�����}�����,> Pbt����� ��//(/:/L/^/�� f/i/�/�/ �/�/GYk�.?@? R?���?�?�?�?�? �?�?OO*O<ONO`O rO�O�O�O�O�O�O�O _�/&__J_\_n_�/ �/??�_�_�__?o �?4oFoXojo|o�o�o �o�o�o�o�o0 BTfx��3_� ������_�_�_ b�t����_��oΏ�� ���(�:�L�^�p� ��������ʟܟ� � �$�6��F�I�j��� ����'�9�K�ŏ� � 2�����h�z������� ¿Կ���
��.�@� R�d�vψϚϬϾ��� ��y����*�<�N��� ӯ����ߺ���?��� c��&�8�J�\�n�� ������������� "�4�F�X�j�|�ߠ� ����������m�ߑ� BTf��v�߮� ���,>P bt������ �//��&/)/J/p/ �/�/+��/ ? ?��H?Z?l?~?�? �?�?�?�?�?�?O O 2ODOVOhOzO�O�O�O �OY/�O�O
__._�/ �/�/�/�_�_�_?�_ C?�_oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\�O� o����M___q_ "�4�F��_V��_���� ��ď֏�����0� B�T�f�x��������� ҟ�����	�*�P� b�t������ί� �e�w�(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� ��9��ϵ�����߁� ������h�zߌ����� #�������
��.�@� R�d�v������� ������*�<���`� O���������-�?�Q� &��6��n� ������� "4FXj|�� ���m���
/0/ B/T/������e�/�/ �/EW??,?>?P? b?t?�?�?�?�?�?�? �?OO(O:OLO^OpO �O/�O�O�O�O�Oa/ s/�/�/H_Z_l_�/�_ ?�_�_�_�_�_o o 2oDoVohozo�o�o�o �o�o�o�o
�O@ /dv��__1_ ���y_��_N�`� r���������̏ޏ�� ��&�8�J�\�n��� ������MƟɟ�� "�4����E����� ��%�7������0� B�T�f�x��������� ҿ�����,�>�P� b�����uϪϼ���A� S�e�w�(�:�L߿�p� 㯔ߦ߸������� � �$�6�H�Z�l�~�� ������������ � �D�V�h�z������ ������Y���}�.@ Rdv����� ��*<N` r��-����� //������%n/�/ �/�/�/�/�/? "?4?F?X?j?|?�?�? �?�?�?�?�?OO0O BO�fOUO�O�O�O!/ 3/E/W/__,_�/P_ �/t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�osO  �o$6HZ�O�O�O ���9_�]_� � 2�D�V�h�z������� ԏ���
��.�@� R�d�v�������П ���gy��N�`� r�������̯ޯ� ��&�8�J�\�n��� ������ȿڿ���� "Ϲ�F�5�j�|ώ�� �%�7�������0� ��T�f�xߊߜ߮��� ��������,�>�P� b�t�����S��� ����(�:��Ͽ��� ������߶�=���  $6HZl~� ������  2DV��fi�� ��G�Y�k���./@/ R/�����/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�? O�&OOJO\OnO� �//�O�O�O_/_ �/4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o3O�o �o�o�o�O�O�O bt��O�_�� ���(�:�L�^�p� ��������ʏ܏� � �$�6��oF�I�j��� ����'9K�� � 2���h�z������� ¯ԯ���
��.�@� R�d�v���������п �y����*�<�N��� ӟ����Ϻ���?��� c��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|�Ϡ� ����������m�ϑ� B�T�f���v��Ϯ��� ������,>P bt������ ���&)Jp ����+���� / /����H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�? �?Y�?�?
OO.O� ����O�O�O/�O C/�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\o�?�o oo�o�o�o�oMO_OqO "4F�OV�O�� �������0� B�T�f�x��������� ҏ����o�	�*�P� b�t��o�o�Ο�� �ew(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ��9�ƿ�����ρ� ������h�zό����� #�������
��.�@� R�d�v߈ߚ߬߾��� ������*�<�ӿ`� O�����-�?�Q� ��&���6���n��� �������������� "4FXj|�� ���m���
0 BT������e��� �E�W�//,/>/P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?�?a s��HOZOlO��O /�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_�_�_�_
oo�?@o /odovo�o�oOO1O �o�oyO�ON` r������� ��&�8�J�\�n��� ������MoƏɏ�� "�4��o�o�oE���� ��%7�����0� B�T�f�x��������� ү�����,�>�P� b�����u�����οA� S�e�w�(�:�LϿ�p� 㟔Ϧϸ������� � �$�6�H�Z�l�~ߐ� �ߴ��������ߓ� � �D�V�h�z����� ������Y���}�.�@� R�d�v����������� ����*<N` r��-���� ����%�n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?�f?U?�?�?�?! 3EWOO,O�PO �tO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_s? o �_$o6oHoZo�?�?�? �o�o�o9O�o]O  2DVhz��� ����
��.�@� R�d�v�o������Џ ��goyo�oN�`� r��o�o����̟ޟ� ��&�8�J�\�n��� ������ȯگ���� "���F�5�j�|���� �%�7������0� ��T�f�xϊϜϮ��� ��������,�>�P� b�t߆ߘߪ߼�S��� ����(�:ﭿ��ѿ ����϶�=��� � �$�6�H�Z�l�~��� ������������  2DV��fi�� ��G�Y�k���.@ R�������� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ?�&??J?\?n?� ��?�?�?_O �4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_3?�_ �_�_�_oo�?�?�? boto�o�?�oO�o�o �o(:L^p ������� � �$�6��_F�I�j��� ����'o9oKo�o� � 2��o�oh�z������� ԟ���
��.�@� R�d�v���������Я �y����*�<�N��� ӏ�������̿?�� c��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|���� ����������m���� B�T�f�ٿv������� ��������,�>�P� b�t������������� ����&)Jp ����+���  ���HZl~� ������/ / 2/D/V/h/z/�/�/�/ �/Y�/�/
??.?� ����?�?�?�? C�?OO*O<ONO`O rO�O�O�O�O�O�O�O __&_8_J_\_�/�_ o_�_�_�_�_M?_?q? "o4oFo�?Vo�?�o�o �o�o�o�o�o0 BTfx���� ����_�	�*�P� b�t��_�_o�oΏ�� �eowo(�:�L�^�p� ��������ʟܟ� � �$�6�H�Z�l�~��� ��9�Ư�������� ������h�z������� #�Կ���
��.�@� R�d�vψϚϬϾ��� ������*�<�ӯ`� O߄ߖߨߺ�-�?�Q� ��&6ｿn�� ������������� "�4�F�X�j�|����� ������m�����
0 BT������e�� �E�W�,>P bt������ �//(/:/L/^/p/ �/�/�/�/�/�/a s��H?Z?l?��? �?�?�?�?�?O O 2ODOVOhOzO�O�O�O �O�O�O�O
__�/@_ /_d_v_�_�_??1? �_�_oy?o�?No`o ro�o�o�o�o�o�o�o &8J\n� ���M_���� "�