��   v��A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@ � &�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	��&USRVI| 1  < `��R*�R��QPRIƍm� t1�PTR�IP�"m�$$C�LASP ��)�a��R��R `\ �SI�	g  �Z�$'�2 �\���R	� ,��d?���aa1`jb�ed`a���a��[`?�  cd�o��
 ��a�o�o �o%7 �o\ n����E�� ��"�4��X�j�|��������ď�)/S�OFTP�@/GE�N�1?curre�nt=menup�age,1422,1ŏ�%�7�ƏT� m��������ǟV�� ���!�3�E�ԟi�{� ������ïR�d���� �/�A�S��w�����𭿿�ѿ�� _TPTX��l�����a` s縄��$/softp�art/genl�ink?help=/md/tp�.dg޿xϊϜϮ� g���������,߻� P�b�t߆ߘߪ�9߻� ������(�:���^��p���������a�`��f�g ($R������6�!�Z��i  ada��c������N��k
������dJ�  ��J�	H����D��4`�~�~��b���`  ���H G?p��K#J�FF��I�:c�B� 1)hR �\��_�� �REG VED�?���whol�emod.htm��	singl��doubt�ripbrows3b�i{ �W�����"/����dev.Es�lo/� 1r,	t�/A�//K/�/ �/?�/5?G?Y?k?}?�?� `�?�?�? �?OO*O<ONO`OjF 2P�?�O�OqO�O�O�O �E�	�?�?_/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoao/' yoso�o�o�o�o�o�o 1CUgy� ������? �2� D�V�h�z������� �O���Ǐُ.�@��O 	_���������П˟ ݟ���%�7�`�[� m���������oկϯ ���!�3�E�W�i�{� ������ÿտ���� �/�A��|ώϠϲ� �����������B� T�#�5ߊߜ�S�e�K� �������,�'�9�K� t�o��������� ����߯1�+�Y�k� }��������������� 1CUgy� �k���� 2 DVhzuߞ� ������ߧ@/;/ M/_/�/�/�/�/�/�/ �/�/??%?7?`?[? m?;��?�?�?�?�?�? �?O!O3OEOWOiO{O �O�O�O�O�O�O�O� 4_F_X_j_|_�_�_�_ �_�_��_o�_�_Bo�Tobj�$UI_T�OPMENU 1�-`�aR� 
d�aQ)�*defaul�t_ ]*le�vel0 *[	G �o�0�o�o��o	rtpio[2�3]�8tpst[1=xY�o�o��=h58e01?_l.png��6?menu5�y�p��q13�z�r�z�t4�{��q��?�f�x� ��������RT�������1�C�҄pr�im=�qpage,1422,1J� ��������˟֏����%�7�I�ؖ^�c?lass,5R����������ϯڔf�13֯��0�B�T�ۓ^�53p�������(ƿؿۓ^�8�� %�7�I�[�ڟϑϣ�������Y�`�a�o ��mΙq�;�mCv�tyN}6Hqmf[�0PN�	��c[1364=w��59=x�q�)�[��tc8�|�r2 ��}Q����w�{�� O������� ��$� o�H�Z�l�~�����Q�c�80������	-`�r�22gy� ��>p���	 -����n����e�w�1���//�*/</7�^�ainedi	�s/�/�/�/��/2�confi�g=single}&^�wintpj� �/??*?<?����r?|!ٙ�gl[55��@�Sߵ?�;Ip�08���076=y�?�5���62,O[I�?	OoO�zl��z�4s�x �O���x� �B�Q�*_ <_N_`_r_�_3��_�_ �_�_�_o�_&o8oJo�\ono�o�o�!;�$d�oub�%oc�13�~�&dual�i38��,4�o�o�o9�o�n�o�ax� �#o������
�%3.=_!g�Q�b8"�z�������\ԏ ���
���+:6��i48,2Q��b]������ ]?ҟ�/� UE߻����s���_���G�u��:���"�f7.�ݣB�Or��4J�\�6G�u7�� ���ÿտ翮��27��)�;�M�_�q�  ��U����������
�!�1�/�A�S� e�wߪ�߭߿����� �߄��+�=�O�a�s� ����������������6
�?�Q�c�u����$��74����������C���6��	TPTX[209�<aAY2+H,���BY1�8t?Ht��(�at0�2��aA0��=�DtvB��O�L_�0��Li�S�=�treevie�w�#X�3��`�381,26�o//A/S/ �w/�/�/�/�/�/`/ �/??+?=?O?�o��
��o%���?�?�?��Ar?>1`��?"2 ��GOYOd?v?�_�.E -��O�O�OxO��@�O 0OC_U_g_��6�OF� '_n_�_�_�_8�_�� �_�S�_Qocouo$vo �o핪o#�oS�o�o 1CUz�os ������
�� y�3�Z�l�~������� �/؏���� �2��� V�h�z�������?� ���
��.�@�ϟd� v���������M���� ��*�<�˯N�r��� ������̿[���� &�8�J�ٿnπϒϤ� ����wo�o�ϭo"߉ '�E�W�i�{ߎߟ߱� ��1�������/�A� S�e�w�9��������� ����e�>�P�b�t� ����'��������� ��:L^p�� �5��� $ �HZl~��1 ����/ /2/� V/h/z/�/�/�/?/�/ �/�/
??.?����d? ߈?�ߍ�?�?�?�? �?OO)O�?5O_OqO �O�O�O�O�O�O��_ &_8_J_\_n_�_�/�_ �_�_�_�_�_�_"o4o FoXojo|oo�o�o�o �o�o�o�o0BT fx����� ���,�>�P�b�t� ����'���Ώ���� ���:�L�^�p����� C?U?ʟy?�UO�O� #�5�G�Y�k�~����� ��ůׯ�����1� C�_z�������¿Կ ��
��.�@�R�d� �ϚϬϾ�����q� ��*�<�N�`���r� �ߨߺ��������� &�8�J�\�n��ߒ�� ��������{���"�4� F�X�j�|�������������������*d?efault؞�*level8�a���Y�w�! �tpst[1]�	�y�tpi�o[23���u�d�,>me�nu7_l.pn5gA^13cp�5x]�[4�u6cp���	//-/ ?/��c/u/�/�/�/�/ L/�/�/??)?;?M?~�"prim=^�page,74,1R?�?�?�?�?�?�"�f6class,13�?OO0OBOTO�?�25ZO�O�O�O�O�O�#�<~O_$_6_0H_Z_]?o218v?�_@�_�_�_�_�O�26�_�o-o?oQocoB�$�UI_USERV?IEW 1�����R 
��jo䒞o�o=m�o�o	-?�o cu���N�� ����o$�6�H�� ��������ˏn��� �%�7�I��m���� ����`�ԟ�X�!� 3�E�W�i�������� ïկx�����/�A�~�*zoomT�ZOOMIN� S�񯺿̿޿�ϥ� &�8�J�\�n�ϒϤ�������<*max�resn�MAXRES���ω�R�d�v� �ߚ�=߾�������� ��*�<�N�`�r�߃� ����������&� 8���\�n�������G� ����������3 A��|����g ��0B�f x���Y��� Q/,/>/P/b//�/ �/�/�/�/q/�/?? (?:?�K?Y?k?�/�? �?�?�?�? O�?$O6O HOZOlOO�O�O�O�O �O�?�O�O	_{OD_V_ h_z_�_/_�_�_�_�_ �_
o�_.o@oRodovo a