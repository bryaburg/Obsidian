��   6�A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	  /GR�P:� $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2� RING,��<$]_d��REL3� 1� N �CLo:o � �AX{ � $PS_�T�I���TIME� �J� _CMYD��"FB�VA >�&CL_OV�� oFRMZ�$DE�DX�$NA� =%�CURL�qW���TCK�%��FMSV>�M_LIF	���'83:c$�-9_09:_��=�%3d6W�� �"�PCCOM,��FB� M�0�oMAL_�ECI��P:!o"DTY�kR_|"�5:#�1E�ND�4��o1� l5M����PL� W ���STA:#TRQ#_M��� KNiF�S� uHYsJ� hGI�JI�JI�D �$��ASS> �����A�����@V�ERSI� �G�  �Z��$S 1�H� ���N ���>_)_b_MV���" ��X���mJ <���:��(_�_t_ �_H_�Yk�Y�A$om�
) �q  �m����#���f�e�4o ro�_7l�o�o�o�o�o��d� ugg@qBq 'w�oooXC|��do��<���=L����3?����@��D� V�h�z�������ԏ0���
�] �E5�pC�-�c��D  2� ������ʟܟ� ��$�6���<��`�r��� ������̯ޯ���&�a|(mZ�i~�i� ����ƿ��ÿ��� π�D�/�h�S�xϞ���$4 1\����I��"If���Iu�P@�]MR�I����ˊ�N%OO�*�N�`E���H@�'I�{q}�B  "��{��!+�����s�2�>@����U�q��-�}�s�y� �2�l�����Qf	6n���j���
�C�[�P�?H!Qg�:�k��� �W���J�ѪN�ER��V��Z�;�^Ѓ:� �u���y���t>>���U�<���,�.�<C�����mAiY>��N-�2�B:w�Q�~ ���B%�@�1LOS)E������|�;� t�_���������,�&� ��J�\�-��Q<a ������r�� ;M���� �"���//f 7/��m/��/|/�/ �//,/�/P/�/3?? W?B?{?�?�/�/?? �?b?�?OOAOSO�? wO�?�?�O(O�O�O�O _ZOlO=_�O�Os_^_ �_�_�_�_ _2_D_V_ 'o�_$o]oHo�o�o�_ �o
oo�oho�o! G�o�o}�o2�� ����`r�� g��d�������ӏ&� ��J�\�-���Q�<�a� ��ڏ쏽��r��ޟ ��;�M�����ğ֟ ��"���ݯȯ��f� 7�����m�译�|��� ǿ�,���P���3�� W�B�{ύ����� ��b�����A�Sߦ�8w���3�,^��ߤ��[��$PLCL_�GRP 1�������� �Dz��?�  ���x�O?r�� ��2��.�A�,�e�P� ��t��������� ��