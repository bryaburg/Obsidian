��   �A��*SYST�EM*��V9.1�0170 9/�18/2019 A 	  ����HAPTIC�_T   8 �$ENABLE�  $BBLNOTEENB=�MAX_ALARMSLIO=��&�ALM-  �$ERRCOD�<' STY;kI}O- X �
�$IOTYP<�$INDEX�T�RG�RSRV1N�VAL=�2��3=�HPCFG�- $ 6�$DEBUG=C�OMP_SWf��$$CLASS ? ���C���f��f8VERS�ION@?  �Z��* </ af��lr�
�r_DF� �2C�(�   �� #�5���C�D�2 ��W���� /./@/R/d/v/�/�/@�/�/�/�/��F�   `�<	"�9G��CG�(�;284`8@9x? �?�?�?�?�?�?�?�d 2?6�
 +O=O OOaOsO�O�O�O�O�O��O�O_�+Uu >
	/K_]S�3U��_�_�_�_�%P_MO#T_	C��R