��   ��A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_  �$$�CLASS  O�����D���DVERSIO�N  ��Z�8LOO�R G��DD<Z$?���q���M,  1 <DYX< [�����D'�i�����iO/a/s/�A/�/�/�/$ ��/�/�/	;�$MN�U>A>"�� � <i#E?  �ı� ę� �ė"0=?O?�5�) g0n2@��4y?�?~�5D�� Ďk0ᗦ0v?�?^9�� �D��0r3�?O@F�A�'"ODOrO�2D�?�/�O���O�O�O�G:��P�ݺu����T:u��g%P�9��:�O=� Y&%P��DɸdC�����QS��P%Pj���;��J:���%P�r�{�껁��Q;|�%P ���
��Ķ���ZUU�I/�_�U��A;6#R:�d��;]�;e���?����h�@�[�y;����?�D�,�5�j��L�Q7NUM  ����a� U{fC2TOOL%?�\ 
;8^�������������]�^���<,!�������n"����C���'c>�Dj�p�I� ��]�׮Q�a? ����.3��4�o;�/��XC����m�a�i4 :f37	o9�iD�mO �_'U;�_� q�����	�� �?�%�Gu�[�4dxc[!j	��