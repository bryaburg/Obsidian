��  	��A��*SYST�EM*��V9.1�0170 9/�18/2019 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP�fBI�IZ@� LRM_REC�O"  � AL]M�"ENB���&sON�!� MDG/� 0 $DEBUG1A�"d�$�3AO� ."��!_�IF� |� E/NABL@C#� �P dC#U5K�!M�A�B �"�
� O�G�f 0CURR�_D1P $Q3LIN�@S1I4$�?���APPINFOE�Q/ �L A� ?1~5/ H� �79EQU�IP 2�0N�AM� ��2_O�VR�$VER�SI� ���~0C�OUPLE,  � $�!PPV1C'ES0�!H1�!"�PR0�2	 � �$SOFT�T�_IDBTOTA/L_EQ� Q1Q@�NOTBU SPI_OINDE]iEXBSCREEN_�4�BSIG�0�OKK@PK_FI�0	$THK�Y�GPANE\D �� DUMMY1�d�D�!�E4�A���ARG1R�
� � $TIT1d ��� +Td+TP� +TP+T5)V6)VU7)V8)V9)W0)W�2W�A+UFW
Q+UZW1
dW1nW1xW 4V�R~�!SBN_CF�![�0$!J� �; 
2�1_CMNT��$FLAGS�]�CHE"$Bb_OPT�2�� �ELLSETUP�  `�0HO��0 PRZ1%ocM�ACRO{bREP	R�hD0D+h@��bl{�eHM MN�yB
1�0UTOB �U�0 �9DEVIC(ST	I�0�� D@13�r�`BEdf"VAL�#ISP_UNI��p_DOv7=yFR_F�@K%D13�x/A�c�C_WA3t��awzOFF_�0N.�DEL�xLF0q8�A�q�b?q�pF�C?�`�A�E�C#��s�ATB�t�1�MyO� �sE � �[M�s��&�RE�V�BIL:�!X�I� �R  �� ODq`^��$NO`M�!QV�l�/�"i��� w����!X�@D�d p E R�D_EV��$F�SSB�&K`KBD�_SE&uAG� G
�2 "_��B�� V�t:5`ˁECY`�a�_EDu � �S C2�}`S�p��4%$l �t$O�P�@EB�qm�_O�KԂUS�1P_C�� m��d\�U �`LACI�!�a����� �:qCOMM� �0$D��Ñt@�pL��O��B BIGALL;OW� (KD2:�2�@VAR)�d!|AB �`BLO@S �� ,K>qA�<`SwpN@M_O]n����CFd XF�0GR�0��M��NFLI���/@U�IRE�84�"� SgWIT=$/0_Nc`]S�"CF_�G�� �A0WARNaMlp�d�`LI��J`NST� CORz-�bFLTR�/TRAT T�`� $ACC�aG�� |L�r$ORI��.&ǧRT�`_SF\gPCHGV0I�Ed�T��DA�Iu�5T���HK�� � �#4aԂN�HDR�B�2�B�J; �C���3��4���5��6��7��8��� 4�z�l@�2� @� TRQ��$�f��ʀ���_Uؖ����`COc <� ������3�2^��LLECA�!�MULTIV4�"��A
2FS٠ILD�8�
1��n@T_%b � 4� STY 2�b(�=4�)2(�P��9Ӱ�� 
7 $��"p��*�=`�L* P�TO���E��EXT���ы��B�ю�22�08��@��%b.'�B s�;�E� �" E�/%ua��L��3s 7�I� Gғ�/A�Ƌ�qM�� � 7��C�! L�0U��� LׯpA²$JO�B6���������IGC�" dǀ������L�-'l��;�Ƨ4�_�M��b# tǀF̝ �CNG�AiBA � Ñ�����/1���� �0����R0��P#p��,}��$��p��t�6q:Q�
2JQ�_RB�qCTJT�YtJ3�D/5C�	�ǧ@��@�  AzO'�n�!% \�0RO��6� �IT}s� NOM_,pn#�cX��ՠTU�@P�S � ��&P���� ǨP�	ѭ��RA�l@n �3�5���
$�TF'%#D3� TD��kpU�1'�q�%aYHr�T1�E ����ң�#Ѥ�%ӢQ�`YNT�"� DB7GDE�!'8�Q�PU���@hֽ��"���AX��"�uTAI&sBUFφ��3!�1�( �װD&J`PIV84'aP�'M�(�M�)6 �&F�'SI�MQS�@NKEE3PAT�nЍ,"��"�!_MC��)G�$��`JB��ĲaDEC[:� [5"����* �I�CHN�S_EMP��$G��7�_��c/��1_FP�TC�6S���5�`��4��q y�V�x�Kx�J�R����SEGFR�Ae�OUaPT_�LIN�?CPVF �A���`�7$+���c�_BNu�DBnrB(	,` +�Ȧ9��A �0��AX0c`5r�D���IX1SIZ\����D��FT�C�Z%Y�ARSa��CD@�IW\%@WX�00@L����0ΌVCRCӥ�sCC w��U%@�X�1խ�2�Mdq�U�1T�XxQ�UDѤ̣�YCk�p����4?`рf��FhEVTFf�F\a_�5F�0�N�ftPX1�h�М)�^Cq�+�VSCAO��A�f�2��(��-հ	��{MGARG���U�F4@Ă��1DWQ�r�0LE	W�!��R�P0Ҹo��l�"R��.� ����ϻ����%ΡR�� HANC��$LG)��a�ǐ��̀:�B�AY���u0RMr��3�s����s4 �xRA���sAZ�0E�B`:�O��FCT�gp��FԠ�R�0D0V ADI��O������������)�)����SpO�[���BMPID�PY �1��AES�7P^c��W��N S�!�qI��/  E�PI,?��40��b@_C�$m�K�� �U0ϑU��1�T#ITq0�V�%97A�."Z_`G2 ��� �!�vNO_HEADE��!~� w�l�0��z�S+��q�R9����43 T���b�5CIRTRH�0�W�XLMt dC��gRJ����!E'RRLX� �4�Q͠OR�B$ᢳ���~{�$RUN_O�p>�P$SYSР4h�͠��U�EV�<W�ǡPXWOyP �=5~�$SKc�"DBT�pTRL
��6̐�P�����7INDI DJ�d��_�`�!������P5L�AS2WAzⰰEE��D!��!R|\��UMMY9���1� |�DBdO���7E��!PR~Q� 
W���-���8� К$f��$Q�L�9$+����P �:Q�ã�PC��;pς�EN5E70Tq<��cþ��RECORj�=�H aO�@78$L��9$Þ"�9���F@t�JA �_D�ʁ� ROS���"SK���rj�ׂ� 1���C�PA��>JBE�TURNA��SMR��U���CR�E�WM8B
0GNA9LJ �"$LA� ���:$P�P;3$Pj�g�<��!b�PC���PDOR@�Q����R�GO_3AW�"�MO���p� �a�DCSSp�STCY��>����0Ls�<�ID���2?�2M�N��OB�>&��j`I� ? P7 $@�RB�Bt��PIM�PO��I_#BY ����TJR&��HNDGj�@ �H�`�1���0{�DSBL=��s�N�0q�,W�(�LS��A��0̶ ,�FB[��FE��@��N�&�)0B? $DO�1�C�pMC�0��I�4���RH��W/ ?(ELE�u
r\�Ǡ(����Cq�$^�q�I�NK)[�UV�LƦ�HA]�QoP$�|#oP#��� D ݬi�MDL �2CΑ5��C���JoR� oR��	��g��	��:�B�SLA5VrElBING ��p�#��&�C�FP�@ P`�p��q�������ou�СO!���!��I!D������W��gNTV�#�VE�$СSKI��`A�C/3	'2IB�1J�f�1����4SAFJ�C'_S}V*�EXCLUs�:��LrONL�0k#�Y���s����HI_yVɀ�RPPLY���R7sH� ~�#_M��b��VRFY_􏳗"Mas$IOj0���&��1IB�$##O���%LSR���%4Ǳ2N�.@a��P-�$,��&AH CNf@�a5N�F3t��G'CHD�s�_�L�LE *�CP��4TǱt�!_X� G���H�TAn���!� ]eNOC
tHlB�pTQоA ~7D��$�I D 9$��6�-:C�!qPCF_\ NLH�LC#��E�@K2�J���q�0x$(B� I� 2_SG�` �K �ΐCUR ~ЛѰ���A#�fЈ��(��H(��FANNUN��j5�CN��@�������YQ��$Z@V֘�EFРI��L �@�`FR��	$TOT�Ч��03�ձ�(5�ǠEM+�NIBK�M6�R��RA���TDAY�LOA�D��䴧R�5���EFF_AXIJ�%N��ڱ�O`=�*��_��QqO2@�`(�6`BcE�Kc�e� Nh Qw1a����A$p&aqP 0�9Q�an� �a�ӯvDiU�Яu�^�CA QjR���n ,�IDLE_PWGsh�e�-�V��V_�`|� ���DIAG_�R� 1$V��SEs�T}�6q� <zǰR���Q�V��@SW�sq��Cp�`�1e� O�1aOHGe�aPPL�IR��B>� �b�ᑠ�:P�r6���x�R��u���e� Q�h 6`,�:uRQDW&�uMSG�6�A��u<arLIFE��BSQ@��"Ns�=r|�Q$q�=rC8�SC�@@��N�YՐ�FLA�3QOV Ј��|��SUPPOn��"��_��E��C_X*����Z�W� ��q�	���XZ_A�Y2�o�CF�T(�)�;uN�9uQ� �vn@��ICTlS =`��CACHC���ؒ`�Et#��y�SU7FFI�����=��b�6��	`DwMSWɕT 8(PKEYIMAGf�TM���SU��BQ�J|g�OCVIE}p��U hBGL�P�?�t@W��0jʔV2@��ST !��YpŤհŤ�PxŤ`ŠEMAI� �=��Q%��1FAULbK�W��<�u�AX�1U�x�pTB>PnXC�R����X��&�0|���LDEBU ����%�T���aYO< $y���S�`v�`IT��BUF�Ȥꗋ�N�!wpSU	B����C�#�z��q�SAV𵲲7p�� Yчp�  VP������~t�_��ֵ�PLɣOT0���cP� M0�v��2s�AX�S]Pb� X��M#$�_Gs�
G�DYN_�q.�PZ <@`D����+��rM�bT�80Fg�%�0DI�2EDT_{���QI[E� GƱxQ&�C������a��ҷQ\�� �� %�T�C_R��IK�rb��B�_�=RM�^��B�D�SPe�B�P� ��I�M���ѥ5B�*pU�y�ހg�`�M�IP`�Bӱq����TH���y��`T�q��HS�~�BSC����`�V�P�J��R�_D^4CONVW!G4�R䍐�֥�Fsq"d0~������qSCr��T�MER�$B�FBgCMP�#A�ET� ]C�FU��D�U��/�o e�]2CaD���g�����NOa1�Q^2B;��U�;��UP�1=�C@�J��1p�u�8�z��P_/H *J�L� �0����>P��#���1 ���Q���Q��a��-�*��7��8��9��s�T����1��1��1��U1��1
1
1
�1,
2:
2����2���2��2��2
2�
2
2,
3:
3R��3����3��3��U3
3
3
3,
94:��EXT-q�Q`�������������t'_��0FDRt/aT��VC0n�pv�D!J�v�REMUp9F��OVMu�j%�As)TROVs)D�T���*MX�,INps)���*qIND� B��
�(	�v���G�� �s� ��|�bqDFf� �RIV�0����GE[ARu�IOYuKc"��N��Q8aW�S�q�|���Z_MCMg��v�1 ߀U@��b y,H�ȱ? �Ar���0rq?�1yE9p�1��Ɽ��9"c`!�P���)pRI�5�ET�UP2_ d ��P��TDDЪa��T��@�1GE����BAC��e T����(ԅ)"�%nS�����IFI�q����@oE�PTrt��FLUI4�f �j�_�{�UR�q۱�����Jਨ�1sV`IW$$�BS��@?x�@J%�C9O?�b�VRT�yPx$SHOUaJP�ASSZ�m����$BG_`MQnMQ���MQ��MQ��FORC��3�CDATA�ag��FU�11�S2�:Ҕ1�A���ah |�� NAV}����@R�_ S����$VISI0�S�C}�SE�07P�eVZ`O�a$a�B�Bx�A�`f$PO�P�I�q�FMR}26%i C" S��bD!6�^fH'O?a?�s?�&I�:uc"_:>FpIT_�A�Tp�M6-??=DGCL=F�uDGDY'xj���DG5��?|��1�M3�jy��i� T�FSJ���k� P��r6�v�$GEX_�q�x�q1����࿂�p3�{5�v�9Gf�6%l �� ��SWٵONA�k�QTLl�h%GR&@f�U��BKU��O1�  �P7`�`K�7���
�:7�M6PLOO��y�SM�`E���A� p_E m ���-!�PTERM��n���AaORIѠ�o���1SM_#в���!p��nq�P�q���q�UP��r� -��!rm�@��)�nr`G.�@pELTX�ҁ�FIo�����0��Ʉ%�o$U;FR)�$>�X������`OT����TqA,�W`��NST��PAT!��PTHJL��E��'��X�ART�b�Yp�����REL���S�HFT��ȑ��_�"PR���� �$��X�q�aE P�Ӵ§SHI'��dU�� O�AYLO���a����@�0-Rȑ�QR��ERV���BC�������`�@�n�@RyC�1R�ASYM���R��WJk��� E �3���B�UB�� ����Yp��P�Ӱ����r�OR�M[c�q��Jds�R7�p�ǐ����a���HAP�TIV�t�2MA 8�������A!��A�欁HO6Pvtu ԰���E6`[`OCQ�|U��1$OP!dFѩ�9S_!$PP�_ T�R���OU,L�ȓe�@Rƕ���o��[De$PWRf 0IM��ĢR_J�`��P�ۓX�UD�2��0�x� v@�$HhE!�ADDR&H��Gʒ-�"���6�RbMaw H�S��	a`Z�nZ���Z���SE�ac��HS�MN�Bx�`B�F"��(�$�O�L�� }�%���R�O�Pa��AND_C���=�¡�Ć�ROU	P��Բ_�0�RU�ձ1�xb0��:�`:� h!;���:���:�yPxb�A`B2��AVED�5��E���Jcy3 $�P��_D�X��-R��PRM_�R^ܲTTP_=�HMawz (H�OBJ`l�[D$&LE�������N`{ � (��@�_�!T��N�qS԰���HKRL��HIT糫�NP��a l�N�%R�F)Sl��Gm��SS� $JQUE?RY_FLA��"�_WEBSOCbG�HW&^�Ma|U�}w�INCPU���QOc�P�& p��%~�%��IO�LNKB} 8�R�I@, $SL\b$INPUT_���$��t�>a MTP SL��Ma~[ q���~���{IO��F_AS�rQ@$Lf@"�fAH�a��o��@a�j��HY'+�A�� UOP�u� ` � I&�"� "s��P����i�"�|�ܱIP_MEan�A� X� IP"����_N
��r���q�I�s�)!��SP0[B��~PBPBG�B� 8�@���A� l�p{�TA��)�A6P㰔`n����`U%�PST&BU�`ID�p��6P�|%z�{%�1#"w"�����5*h$I$| N��(�`�%�IRCA�_CN�  � ��@�� CY��EA
1a<g��'7��C��=�~#x�DAYy_� (NTVA�E�� k7��w#k7SCA��k7CLq�!-Q��"`�A��/�$�,�%�5N_T�C�B� �"Y1�@���P`�A��� {!��_8�Q 2� �$!iA�A�� $RF�R �LAB��pA�`vGU�NI�dC̀IT!Yb$!&�"R��
Pژs��CUI�UR�L�P�$A��EN�?�ۡ�Q����T��T;_UA2 �J �QM��$R"�J�@" Ra$P�`A��2.QJ��9RFL�pA0�x`
MS5s
�UJ]RIe� �� F�p�q�P��yRD�3$�J7��RJ8�Y7��p^2�R�W7uF�P8��Y�QAPHIBp�Q�S�WD�pJ7Jy8ڢ`L_KE�@�  �KG L}M�! � <�0�XR�  3WATCH_VA�Ѱ��A��FIEL��y��0(b�u� �`��V��V��aCT�@�f��LDM� �x4��_M��ΡD<�1Q�LNTK����'COO���fNF��f!Ta�`����JvP��(�����LG�d��� !�)LG_�SIZH�9�[uMRXYw� ZvFDexIYx pxl�gv|x��ZvWpf� `s�vop�v� �v�p�v����v�n�P�_��_CM��#�Lg+�'�AF$�1�K�Wp��(Vqc�bqp�opp�� p��p|�Io����p0p��pp�WpRSK`אo  (2�LN�Qj���U��DE6�E�`��A����԰�L���DAU"�E�A��G 6�8�.�GH�7�dQ� BOOO���� C
�IaT��l�/RE* ���SCRX��D�����"�MARGI ��з���U�ᒍ��S.��W������JGM�MNC�H���FNb�K@��@>�UFL���L��FWDL�HL��STPL�VL��@L�s�L�RS��H��h��C����A������U��`�򗈃��`2S�G0�	�POW��������,�6�!N�EX.�TUI>�I�pC 0�q.�ֳ�ֳ<��A���o���������N�����ANA�+tA�VAI�P�Ա3�eD�CS\0b�R�p�R�O�X�Od�SA3��o�S{�֘IGNpp�0�sp=��`*A[�DEV��LL�aZ��#Cpi��`�!Tr�$fw��H 49r��A� ����0b  �ѭ�S1J�2J�3�J�炈�S�Cp� �@�p)t}��~|%�����r����Q��ST�[R9�Yr�� /�$E��C�ۘP�����	�B��Bq� L �p.���e������j�X���_ � �������3����� �MC���� �� CLDP|[�eTRQLI�AV���FL!��lQ���1Dwa����LD8������ORGQ����RESERV (M�4M�?��lS� ��`�����F��SV����TR	1������RCLMC���M�_���J ��`M�DBG�Q�5`�1sMA�dU0FC�U��T8�r%E�P���MFRQLߙ � KyHR/S_RU�b�DyA0$�FREQ6��u�$�YwOVEARj �s���~VPU�7EFI� %G�Dp3u��[z�� \P���T$U��B3?�`�1PSI�9P�	��`��D"��U|� %?( 	}��MISCkU� d,����RQ7R	 p�U07P�鱎AX��b#`��EXCE�S�BM�cM)@oQ�²`u�d��eSC>�� � HA�_I@>0+��s��K�D��d%B_^�`FLICB�B��QUIRE �pu+QO�+���Ld�M�E� ��{�� �b�c��WND�g0pP!����Lx 3D;�
�INAUT��
�&p�P8��Nr�q��!����!PSTLoQ�� 4�0LOC��R�I�@��EX�6ANqG*r.aODA]��qrBzPbMF�b�u���c⽰m�8�5�$SUPi���FX1PIGG� � ��`c��q�� c�
�c�@���5I�� EH��TF5 t�0�CTIl`C�Q!�pM!Pn� t�0MD�AIB�)�FX��D���GqH�0�Q�DDIA�Q�C4PW��D0ѧ��ED@�)OjS��pP�� �CUppV�	P��.���0ؑ_ � �{Еӿ3L 4r��p|XP|^hr����PP{XKE�T`e�-$BW�oV���ND2��Pc�Q2_{TXl�XTRAX�4�R���� LO:��1��d" f��CR.f&c�RR2>h�� -a��A�� d$CA�LI��uGF�jg2�F�RINb�nc<$Rx`SW0���c��wABC�8D_J�P�{!.�A_J3�f
��b1SP� P.P��d�m3�mHQ9�.B#uJ��3un��O���IM��MCSKP ��bt7�?�btJA�M�Qb|�uyu�u�w�0_cAZ��/q�qEL��<.r��OCMP�3N��RTE�s e11�0pe�1����: �Z�SMGՠ�@v��JG��SCL��5SPH_��M���f���.u`RTEIR�`nc�k`_E�
��b Aؐ��M��sDI�qQ�23UdrkDF!�āLWʈ7VEL��INx���_BLX�.��Yq�/J�����1PIN���]`�CR9�ْ�TR8�6�_T �@F�a���j�^�"�k����+`DH��P\a���$Vw`3_����$=��~&�$���Sah�H? �$BEL�pm���_ACCE�� �	����IRC_4��q@�NT��O$PS���L!��0M���9�.��1G�@/��Q���$���3S�T@�_G�ؒ������8�_MG}DDء��~FW��@����$���DE�PoPABN[�ROg�EEˢK�B����qK�� �!�$US�E_v`�P$ CTER�Y4�ꐪ� ��YNgA鰢�Rp�AB��M:NQ=�ҠO�v�ϴINC(T�1������Yq�ENC��L�A.K���H�IN��IS�8ť@O��NT��NT231_Ȃ~f�LOـ~|�� I� #��΀# $ ��h��#"CQ�M�MOSIݡ<"[P����MPERCH  �ó�� �Ǚ1�� lA����lA�w�r����$��PsAS�E�L��Ps�7'OwN�@�ʄ֟�T3RK��R�AY"c?� !��S��ոӔ0�v!��P MOM鲎" C�HP$�jg�ӆ��g�T`DUXp��S_�BCKLSH_C M�F�: �ƴ ��-e���o깱�uCLAL�MJ�@�Њ���CH�Kep�@�TGLRT�Yp@�S8ėE5�A_��3��_UM3��C�3�Z�� LMT�`_LG��s%��A0�E*�K�=�)�@�F�@�`p9NҌ�)�PC���)�H@� ܥ��CMqC�U��CN_�b1N�S��;sSF���V���A.ǃ���M�/n��CAT��SH�3 �b� ���/�/�eT��i�٠PA���_	P����_fpZ�����0eq�����JG�0���ӀOG����TORQU~��e���� �`e"�� �B_W� ���ّaʓ`Г`UIhIvIГF�0`S:r�Iq�VC�0!%�1�ڠ��q�JRK�!"&�<PDBX�MtS<PM�0_DLʑ_�GR�Vg`$ʓ`$ГA!H�_%c?#���*COS�+�p�(LN# �+� �$ʐ�)=��)��*�,İ<%Z� ��A!MY��!:8�"�Q�+[9TH�ET0��NK23�Г�2ē� CB�6C5BēCz`AS�A�2`��1ʓ�1�6SBʓ��2�5GTSkqZ�C��a���&�J�#$DU��h�6Bjb���EG�Q%�_��xN	EhtP`I� �������y1A}5�E�G�%�(�!LPH�%�B^ńBS��C�%�C�%�B6P!SZ(6�@V�HV�HT���LV�JV�KV
[UV[V&[V4[VBYH�H�F�R�Md�X�KUH
[H[H&[H4[UHBYO�LO�HOsi��NO�JO�KO
[O�[O&[O4[O(6F��B�1y�%t�GSP�BALANCE_lJ16sLE�0H_}5SP>��&^r�&^r�&PFULCbx�rqw؉r�%K�1��UT�O_����T1T2�y
�2N���V��t�M��ыpi@Z��	�T�u�O���QINSsEG���REV����G�DIF��p�1٫U���1���OBK���j#�2,V���~I$LCHWAR4�摲AB��$MECH�1J0��ǁ��AX��Po����G���p� 
�?�0�7ROB��CRM�#����@�C�_�T� � x $�WEIGH��w �$�C\�� I����I9Fv��LAG����qS��:���BIL��cOD�Ы�s�ST�"s�P:���t��N C�L��P�
������  2���x�D�EBU��L|�Ē�5@MMY9C�9�N8�$�w $D|� ��$�� l1 �  �DO_:�AK�� <_�ޖ�p��$���@B����NJÁ��_���� ˒O�� ��� %�T�7�?��TL��F�TgICK����T1N�%֣=�ߠN���pu���R\ఱ��񥩂���U�PROMP��E~�B $IR"ற��8�X�w�MAI�F ���Q�_���O�X���°RU CO�D�FU����ID�_����8�2�>pG_�SUFF� h����X��DO��0/�������GR���� Ѵ�ݴ��赩���-�ѴU�퐱_�H�_�FI�9G�OR�D�� R��36�s�H®�N�$ZD�T��M�ˑX��4{ *W�L_NA���ߠ���DEF_I �ȡ��������𦿔`��������ISm@@# m�|@�0�����D6�4���D�p(?�f��DO@pl�LOCKE�˳�`��2�Ѳ˰UMе ��Ѵ��Ѵ��Ѵ>�ݲ ��ܵ��ݴ�ݲ��2� 2�賴��赡���� �9�w�͸��P}� ���,т@F�W�ر�����TE��Y�� ��LOOMB_����0s�wVIS� ITYs��A�O��A_FR1I�s�~�SI,��BnaRܠ7��7�3��
s�W�W�Q �% 9_���EAS{��@��| x�W�8�45��55�6|�ORMU�LA_I��G��ǵ h 
�7��COEFF_O á&�)á�0Go{�S��5�CA�p:�L��ˑGRm@ � �� $���rv�X��TM�ד��ɢ��,��ERI�T�Ԑ�n퐳  �rLL�:p�S�A_SVk��$��퐴.0����� �SETU,�MEAG����t��ˑH�L�� � (� ���lقl��w��ߠ�ќ�	}�]d������y�G�xг[@��Nk�REC[�q���SK_Apy� �P_�1_USER��q�2$��*4 �qVEL� ��-"!%���Iz�B��MT��C�FG��  ��]�OςNORE�J���l"�OPWO}R�@ �,B��SYSBU�P�S�OP�!��T�*Uğ+X�P��K"�%PA` q�#˂�OP�U���!}����� OIMAGz�� fd�IM� 5IN����"3RGOVRDfP�#	 �!P� 3 ��|@g�l�i5ЂL��B�T:BlPMC_E(���!�N�`M�2���1� 	�H1S�L|p�� �R�O�VSL�S��DE�X\���5a@��8_ H0�7�I0�3��3GH�4CC����5CA�GI0_ZERl!��2:�� @ 4_C�O��RI����
�Fg��I�A�AQZ�9EGA�� H_�̀�ÐATUSk,�C[_T31DX�FB�  �F�ApV���C���� Dc�� �2�B�P�-��AM�- �r1XE@�@x9RMRTvC�}@�`��@UP�H�&�P!X;�V�1�3�7R���PGY%�� $SUB�A�E��A��CJMPWAIT��PC�ULOWςF�ʡM��ЁRCVF�_��ς�QRE`F40���CF@RLς��<gIGNR_PL^�CDBTBÐP*�FЁBW�2dt U���1eIG�!!��qҀTgNLN0f�bRT{3�NO�N!��3PE�ED�P�3HADO�WÐ΃t ERVE`�3�d�2�Q��SP�p � L_�瀼��`1�tUNq��[p2�QRTPNCLYw����AP!PH_PK�TZ#�b"RETGRIE�Cx"�"r�WpD�FI_r� �xR�Zp�t 2�d �DBGLV@cLOGSIZ܁�Zpa�Um��tD�c�`_T�XτM��C�B�E�M�}R�s��ˆCH�ECK~`� �PL �� 0@vx9�gALE�Qx�PA��0����SrIP�b��
AR�r��N�=����@O��b��AT@��xc��v�pل���1sUX� ZBjQPL���Z$� $d!��S�WITCH�rE�W�O��A�R�LL�B��� $�BA�DvӞBAAM�@.�C=��A,�#J5�`N!Y�6_��_KNOWO�u�L0�U�AD/�c 
pD� ��PAYLOAq9ී_�A���!���Z��L�Aj��L�CL_�  !@4��S�?!�]2�F�C� ��p�� I��R� ��W�@P��B��� _J@r~�_�J�� !SPTANDq�������~!���PL�AL_ )��
pA�B�1���C�D��E��J�3��Ŧ� T P�DCK�0)ҞCO�MH�PHգ�BE0.��կ��X|a>�0 � ��`��WD_1��2�DMAR@Q��������:P_RTIA4ù5ù6�MOM��ϳ��ܳ��V B`AD�ϳ�ܳ��PUB�0R��@�ܳ@�:�+������ L$PI�4�at�!�ɨ=Aܙ��I��I��I �à���\��ơQ�ƬQ$RO�c��E�cHIG��ce�d 4��de9`.`4�j�C��9aR�9aeSAMP HP=���4ק�eN��� &��� ��!" �ԡP���`���ٔ�!"�R��ȴ�Տ�m���IN5����<�X�3�b�>�~�U�~��GAM�M*�S�A���qGET!�FIO��c�>"M
WIBF�bIl��d�$HI���AH�@!"�E;� �A�=�.�LW�[�R�=�@�.�X֚`ǡCheGCHKV0�@�
�#I_�Й�>"1�r� v�$������1���ţ� �$�� �1���IRCH�_D#��P$d�L�E;!!�At^�< ʾ�`MSWFL3dMn��SCR�X752 �p��O����F�ϰ`���	�`�k�SV#�w�P�pCUR�#f�pSAA�n4A�NOb�C�A�c� A��r�ȟڟ�Ȯ�`���������DO�aA���q���
�.ؚ"�>�^�j�?';%��� ��bLS r�� � ��YL��r�$����p�%�r�'@`�@	�"�#r�(0� @aN7QM_Wp�"�"`��#��s!MG`�+��'ġd�4���5�Rrl�M2wB� ��q�� �4$WQ0�5ANGLa�Q0:�O2�A�O2H�O2�X`;�N�o������sw�XGpO�I�v�Z�5l�`r��[ ���OM� �����ư�pg�*�j�b�_�R� | �HN﹛Fܳ�F:� NȺ�G�F����p(B�p�D�P���PMON_�QU�� � 8�:�QCOU:�Q�TH|`HO�"FPH�YS��EST�FPU�E1P7UpO�T� � gpP`�bRU�N_TO�#�`O!�� P���U!e�#INDE�sc�G�RA� ܀� 2� N�E_NO�T�UITxj �QsPINFO��er�[a�"�L1O�Ib� (��SLEQ%�.a�.`�V�0�OS��p�� 4�:�ENAB}2�PPTION���d�g��dbcGCF�q� �@:�J0v�R���R�hhq�o�d���EDIT� ���p�0KE�&�$�E�,�NUwxAUT<]uCOPYE�!�(6|�iM�N@pD{^��PRUTq2 Gr�N�`OU �$G��R�t'RRGADJZq�y�X_� I\P�0�v�0�vW�xP�x�� �v=ӻpBbN��_�CYC}2i�RG�NSge� w�LG�O���NYQ_FREQW�W���\����SL򐞂T��q���&�CRE��QS��IF���SNA���%��_GjSTA�TU�@j�WMAI�L�Ҁ�IuATLA�ST��.�ELE�Mka� ���vgFEASIxa?"���  � �&�JE��b!���I�P��S��IQPy&z�AB�a�E�PAЁV���~�����X�U�_�!�V��ǖRMS_TRt�v�g ���3^�Bb �Ɣ XM00��3݊@	Q�? 2� d�4 R�7���6��.0 �!p��b���nDOU�S2bN�c0�PRd l`=�5bGRID�Q�coBARS%�TYycεrOTO
�q� �Q_��!�pݢ���O�0hd� � � �@POR�S���.�SRV��)&��DI_T��?�R�Ј\��\�4Z�� \�6JZ�7Z�8>�o!F���ka�~P$VALAU��47�vArPF4��� !teX�Qb���1�`AN3��́Rpa�5�TO�TAL�Ӱ1A�PW�I�I��W�REGENU�j��CXӘ�Sa�Q�,PTR��W�U�C_S7��j��cV�q�d�¢b��E샩�KQp4��R,p�V_HƠ�DA,C���S_Yhe�2m�S� AR,@�2� �rIG_CSE�������_�P���C_Ѧ$CMP,p7��DEtKБ҅I��Z��\�Ba��E�NHANC2Q� p$�ve̂ ��GINT=�g�0F�S��1MASKȃĐOVRQSP#P��H@��@vầ�V�e ���pb�V���Ѧ�PSL)GT�ka�`=n��02?�H�S�"�����U�2��TE�0İ����o���Jb�]}�IL_M`|��w���@TQ,P���Q͐��"V2�CF@�P_�VJ�Ma�[V1`�V1n�2}�U2n�3}�3n�4}�4n�#��!"#�`����!"IN	VIB�<0:�' !.2*2�63*364*4�6p:��Np��T $MC_F,OPd$ LBN��5�MnI�Ӳ~�� �@5B��� KE�EP_HNADD"�!����	C�1��Aݡ���O%Q��zp�2 ��REM%G� �J�afU��eHP�WD  �S�BM���COLL�AB.4���3����`IT3��0UrNO5AFCALt2��47� ,7`FLz0���$SYN� ,M��@Co��V�UP_�DLYq�~RDE�LA= H�ɂYPA�D,A�QSKI�PS5� ���POƟ0NT�!g P_ �P�R�'�P�2g��'�� �)�a�)s��*���*����*���*���*���*9��q�RAhd� X�J�'���MB3NFGLIC�S[0T�US�<���WNO_H[ D�Hq�2IT�r<0_�PA�PG�� ����UҐW�`�6M�>��NGRLT= �Q��q��������1�Tc_J�!�6BbAP���WEIGH�SJ43CHxP�4OR��4�$�OO+���d��6J	���AaA��nCIHcOB`�`���J2s0*q�pcX��TV��A �Q5��A�p��A�Q�?���RDC��W� �
pR�cR0P9�"R���JIR�B9��RGE�`c��C��F�LG7�PH�d9�SsPC�S�UM_�@>��2TH2N��_@��A 1� ��s0ݡ4� � �D����I��2_P�d2�SS����]�L/10_C{��1�Tn�� ��p$�P 2�Y��C�;�� a�D��aZ��Q�C7cp���hқ� �V��МP� P��DE�SIG�RV�VL1b�Y1�VTcg10a�_DS���2EFvOp11q� l� `��!��ATCp�t��_��bIND�����aOp9��b�2H�OMEr �e2�b��o�o�o	-*��d3�b�Pbt���� �@�b4�b������'�^?p�$$Ch�SBPO���ā773 ��	�SI"��π�Z��$AAVM_WR�K 2 ą� 0  G�5ˁ�%��.H� H�	k�\��7ŀ�m�������[�Νڟj����'��/��BS�`�A 1��� <�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ� ����������
��.�@@�R�d�v��?�C( �AXLMTBP����X�  d��IN�����PREoPEb������_C_��wO  �� c�|�� �ID ?ą�� 8�d�^� p����������������9�-a���J��U�Pb��4  ~�IOCNV_lP�� ȴ�P}�0��pT�>�V@�  1 �P $�畑���ŀ?�L��  $6HZl~�� �����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4oFoXojo|o�o�o�o �o�o�o�o0B Tfx����� ����,�>�P�b� t���������Ώ��� ��(�:�L�^�p��� ������ʟܟ� �� $�6�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿�Կ潝�LARMRECOV M������LMDG K-� L>�?_IF ����d  YST-0�34 HOLD �signal f�rom SOP/�UOP is l�ost ide �Clear,G1�,A1) 11 ���executed VPL�Á�������!�3�W�, 
�<h���8MAIN� ��LINE 2�7��AUTO R�UNNING��W�ORLDo�����$��� _PLAS�TI��ALLET_LEFT K���$����RNG�TOL  �	? A   Y�k����PPINFO H� Gƞ��8����}�  T��� �-���-��Q�;�M����q������������+�1CUg y������3��PPLICATI�ON ?������H�andlingT�ool�� 
V�9.10P/23�z��
1667�7557H745�8918\162�64H=O7D�F1C���Non}e�FRA�� 0��_A�CTIVE�  �R�  #��M�OD ]�P�%CHGAPONL?/�c�V OUPLEDw 1p�� � �/�/�/
+CURE�Q 1	p�  T*�)�,�,	?$5 94.��/??+?=?�O?a?�?�?.���"�%�4�H�%�"�:HTTHKY�?�?�?�?�? 4OFOXOjO|O�O�O�O _�O�O�O__0_B_ T_f_x_�_�_�_o�_ �_�_oo,o>oPobo to�o�o�o�o�o�o (:L^p� �� ������ $�6�H�Z�l�~����� ��Ə؏��� �2� D�V�h�z������� ԟ��
��.�@�R� d�v���������Я�  ���*�<�N�`�r� ����𿺿̿޿��� �&�8�J�\�nπϒ� �϶�����������%�TOC�/1#DO_CLEAN`/$���NM  H� �/����	��-��.DSPDRYR��&%HI= ��@�ߙ� �����������)��;�M�_�q�(MAX@~�7��o'��X~����"�"PLUG�G~ ׋#/%PRC*P�B������z����O��Y�k�SEGFW K5GR���߀�����LLAPv��35GY k}��������/R#TOTAL�����R#USENU
v �+ d�h/�� �RGDISPMM�CU ��C]��@I@k�$Ot���a�#_STRING� 1
O+
�kMH S*
�!�_ITEM1�&  n-
??.?@?R? d?v?�?�?�?�?�?�?��?OO*O<ONO`O�I/O SIG�NAL�%Tr�yout Mod�e�%Inp�@S�imulated��!Out�L�OVERRs� =� 100�"In� cycl�E�!�Prog Abo�r�C�!�DSta�tus�#	Hea�rtbeat�'MH Faul0W9SAlerCYsOa_ s_�_�_�_�_�_�_�_o z��+z��/ oTofoxo�o�o�o�o �o�o�o,>P�bt��oWOR U �+�qDo��
�� .�@�R�d�v������� ��Џ����*�<�N�PO�+$Qt��{ ]�������͟ߟ�� �'�9�K�]�o����������ɯۯ�o�DEVw�����?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ�>��PALT0m�� ���������,�>� P�b�t߆ߘߪ߼����������(��GRI���+`���:��� �����������*� <�N�`�r�����������N�F R0mx��� ,>Pbt��� ����(:�L^p��PREG �Ω����/ /*/</N/`/r/�/�/ �/�/�/�/�/??vM��$ARG_�pD ?	���W1��  �	$vF	[�k8]k7�vG�9J0S�BN_CONFIQG�@W;�A�B�1��1CII_SAVE  vD�1�3J0�TCELLSET�UP W:%  OME_IOvM�vL%MOV_H8@$O*OREPuO�@:UTOBACK��1W9�2FRwA:\� �O,��0'`P��H�� �K�0 �18/07/�10 22:%P18��8�6_H_u_l_�L���_�_�_�_�_oo���_DoVo hozo�o�o)o�o�o�o �o
.�oRdv ���7����p�*�<� �  �A�_�C_\ATBC�KCTL.TMP DATE.D�����������ˏ�CIN�I���E�6�CMESSAG�0��1_0��3�1��ODE_D�@�6�$�O�,�ޒCPAUS�� !��W; , 	���0�%y ���vϾ	���8�]��n @�*ݖ,		 ��W5��Ɨ���П� ���@�*�d�N�`��������̩_�i�TSK  o��A�1��J�UPDT#��d�9�Z�XWZD_E�NB脸:B�STAp�W19�I1XIS�0?UNT 2W5�1��0� 	�@��
��� /��O نn�Y�� �Ȗ���IB Vg �s  ZH ?Q� #������	Ϥ���� gF���B ?u�������� �D��3쿸u�?;��MET 2���3 P��I!���H���H��>wFd�H����I�}�ƶ@��Zx?��e?�c��=M�7?�@4�����SCRDCFG �1W5�A 	��5�2m�A�S�e� w߉ߛ��O�U�9.� �����!�3�E��i� �ߍ���������N���B7�AGR��-�M��&�^�NA>@V;	��D#�_ED�1��� 
 �%{-d�EDT-�0RJ���� ����(�B����2�_��\��D ����29�QKPALLET�j�OP_VERI{FYp  =d0 ��b�,I\V	3QK�`R���.@��&���4� A/ew�e/��T/���5�//�/1/ w�/1?x/�/ ?�/��6i?�/�?�/w�?�? D?V?�?z?��75O�? �O�?w^O�OO"O�O�FO��8_��N_��� x*_�_�O�O�__��!9�_=_oa_�x�_�ao�_�_Po�_��CR 8pO�o�o�M�o+ro��o�o&�s�NO_�DEL2�$�GE_�UNUSE0�"�I}G� OW 1V��   (*SYSTEM*��	$SERV_�GRj���pi�RE�G�u$���pN�UM�8�&�PM�U�p�LAY|���PM� |�g�CYC10r~ⅎo�s���ULS���l����i��sL�����BOXORI��CUR_�&��PMCNVa���10��M�T4D�LѰߏ�	*PR�OGRA�tP�G_MIs�����AQL}�������Bڟ��~$FLUI_RESU������C|C`�r����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�FπX�j�|ώϠ�x&�L�AL_OUT ��{E�WD_A�BOR����IT�R_RTN  r��=�
�NON��3� �xCE_R�IA_I�p5��~�A�h�FCFGG V�~�u����_PA��GP 1]������������C�  �>�@�@�@പ@�@��@��@���@��@��@��  �D��D|�|��8�S��@�@���@��@��|���D/� D|� ���p+D3��=|�F��j�DY��?��h�H=E`pONFIU��n��G_P-�1�� }uV�8�J�\��n�����������KP7AUS�1�~�{ �� �	�����I��jS���������x���� �Ϻ�0�Z@j �v������� DVh�M*�N�FO 1�}�� � 	�����Ћ�������Yr���9���¤@`���g�3i D����?�qC2����޿�����B_���h�OƋ��ߧ�!LL�ECT_��y� �9'EN}�5���U"!NDEA#�I'�s>r1234567890�'�9b�q�ҧ/�&.c
 	H��.c)�/?�l�/ ?^?;?M?�?q?�? �?�?�?�?�?6OOO %O~OIO[OmO�O�O�O �O_�O�O�OV_!_3_`E_�_�ͅ$�q2I+� ��X+�"IO # �)U!.g4�o�.o@oRo�WTR��2%!�](��i
{_`n���"�]�j��]&_WMOR�R#�� ?�? -B����u �y+O=s�{��b���Q$�m,��? ����W��q��K�tyѕ��P"&I/�� ���.�@�t�
�r�(/'���e�i@���\|��c ��a�h�PDB�p(�̉Tcpmidbg����1�*�:�^��p��]�(����^���l�o���K��6m��Ɵmgڟ3�����f"�{�<���Pud1:��ɯ�j~�DEF '4�c)��cّbuf.txtԯ"�կ.��_MC�c)���SQdg�H��d*V����|��x�A�C� �B�!�C9C�aC�C�%)C3�C�-��D�n��D���D:��D�x'D�pj�ESAo�F;��F��F��iE���F�� Gb�7�kr S zD��w,�\rЪ��cĽ���`�Z�c�`x���۱��Cf@�1�D4�\�D��E�H��D��D{�F���3ES�F�I3���F��E��}E{�H�F{��G�����  �>�3��C�r��n8�ѧ���5��ᧁ�cr��A�q7�=L��<#��ea��X����@�RSMOFS�T %�X��P�_T1w�DE -����a;���;�Q�s�m�?����<�M<�T�EST�+��R�C"./vC��A��7����?ї�B0�������C����s���:d��b*[�I�#/e�?��r�0�m�$r�RT_~�PROG ���m�%3�S�X��PNU?SER  r%���f�KEY_TBL�  ����	
��� !"#�$%&'()*+�,-./�':;<=>?@ABC��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������-��������������������������������������������������������������Q'�L�CKq�m�h�q�ST�AT�Y�_AUT�O_DOo&l���INDj$�8!R(����"-24�!# STO�  �TRL)�LETE�o'{_SCRE�EN �j�kcsc"UlMMENU 11� <B�A�	/X� �/G/��$/J/�/Z/ l/�/�/�/�/�/�/�/ 7?? ?m?D?V?�?z? �?�?�?�?�?!O�?
O WO.O@OfO�OvO�O�O �O�O_�O�O_S_*_ <_�_`_r_�_�_�_�_ o�_�_=oo&osoJo \o�o�o�o�o�o�o�o '�o6oFX� |�����#�� �Y�0�B���f�x����׏��������_M�ANUALp�ZCD��2�ل��R���gߗ�?|(��g�L�@�3F� Bȗ�7�z��7�0��$�DBCORIG���	�_ERRL&/�4V����>��P�b� �NUM�LI*�Wg�m�
��PXWORK 15V�-�¯ԯ����
�[�DBTB_�� 6���b��t���DB_AW�AY��GCP� m�= �^�_AL*��^��Yo�m�&`�� 17��� , 
����e�(�v������ݾ�#�_MI��l�@@�4�ONT�IM��m���Tƪ�
����MOT�NENDu���RECORD 1=9�� �DF�A����C�k�D�I�A�D�C���(B@?UB�@�A�r���!Є�Ĕ
�EXECUTIN�GR�&�8�J�#�G�O��l�W߀fߣ�m� ��������_���� ��\�n�����%� ��I����"�4���X� C�����������E� ����{�0��Tfx %��A� ��P�t�� ���=�a/� :/L/^/p/��//�/ '/�/�/ ??�/6?�/ Z?�/~?�?�?�?#?�? G?�?k? O2ODOVO�? zO�?sOO�O�O�O�O�gO+�TOLERE�NCk�Bȴ�y�L����CSS_C�NSTCY 2>J���a�_���l_ z_�_�_�_�_�_�_�_ 
oo.oDoRodovo�o�o�o�oGTDEVI�CE 2?W[ F�#5GYk�}����#�HSHNDGD @W[Ƨ�Cz�z��JQLS 2A�m�G�Y��k�}��������IRPARAM BY��k�v�5��RBT �2D��8�<<ذ C;P���ª  �;P�Q��@W���E�?�d
�Q�HZ�Ԑ�\^���@������M�+C�J��8P V�͐0ŌU��;�B�J�6U�ŅD�@����;�@��h��\�X�ńc�� ņ���Z�l�~����� ���د�7�� �2��ŅC�,�D
�D�0N�� 	��9�M<A�+�A���,A���A�?�A�U2Ŋ��YCs���B���4δ��Ō���|%Bw�q�B�0NB���QB�>_C�񹴿ƿؿ����? ��� gp� ~�H�ō-�O�a� ��I�wωϛϭϿ�� ����B��+�=�O�a� s��ߗߩ��������� ��'�t�K�]��� 7�������
���.�� R�=�v���cϑ���� ��������<% 7�[m���� ���8!nE W�{���g�/ �4/F/1/j/U/�/y/ �/������/��/�/ B??+?x?O?a?s?�? �?�?�?�?�?,OOO 'O9OKO]O�O�O�O�O �O�O�O(_�/L_7_p_ [_�_�_�_�_�_�_�/ �O	_6o�Oo1oCoUo go�o�o�o�o�o�o�o �o	h?Q�u �������� R�d��_��s�����Џ �����*�o3�E� r�I�[��������� ǟٟ&����\�3�E� W���{���گ��ï� ����X�/�A���	� ��Ŀ���ӿ���0� �T�f�A�o����υ� ���ϻ��������� b�9�Kߘ�o߁ߓߥ� ���������L�#�5� G�Y�k�}���E����� ��$��H�3�l�W��� ��}ϫ�������  ��	V-?Qcu ����
�� );�_q�� ��/��*//N/9/�K/�/o/�/�/�/���$DCSS_SL�AVE E�����!�~�*_4D  �.~3CFG F�%�3�dM�C:\� L%04d.CSV�/�{?�  ��A �3CH�0z��/g>�?��?�  �g6���1O�9A� J#(C�;g4��0��7,4RC_OUT� G�+OB�/_�C_FSI ?~�) :K g6�O�O�O�O�O__ F_A_S_e_�_�_�_�_ �_�_�_�_oo+o=o foaoso�o�o�o�o�o �o�o>9K] �������� ��#�5�^�Y�k�}� ������ŏ����� 6�1�C�U�~�y����� Ɵ��ӟ��	��-� V�Q�c�u��������� ����.�)�;�M� v�q���������˿ݿ ���%�N�I�[�m� �ϑϣϵ��������� &�!�3�E�n�i�{ߍ� �߱����������� F�A�S�e����� ����������+�=� f�a�s����������� ����>9K] �������� #5^Yk} �������/ 6/1/C/U/~/y/�/�/ �/�/�/�/?	??-? V?Q?c?u?�?�?�?�? �?�?�?O.O)O;OMO vOqO�O�O�O�O�O�O ___%_N_I_[_m_ �_�_�_�_�_�_�_�_ &o!o3oEonoio{o�o �o�o�o�o�o�o FASe���� ������+�=� f�a�s���������͏ �����>�9�K�]� ��������Οɟ۟� ��#�5�^�Y�k�}� ������ů����� 6�1�C�U�~�y����� ƿ��ӿ��	��-� V�Q�c�uϞϙϫϽ� �������.�)�;�M� v�q߃ߕ߾߹����������$DCS�_C_FSO ?����?� P � �\��������� ������"�4�]�X� j�|������������� ��50BT}x ������ ,UPbt�� �����/-/(/ :/L/u/p/�/�/�/�/ �/�/? ??$?M?H? Z?l?�?�?�?�?�?�? �?�?%O O2ODOmOhO zO�O�O�O�O�O�O�O 
__E_@_R_d_�_�_|�_%�C_RPI<�N�_�_"oo�_;���_.owo�o�o(�SL�_@l`�o�c�o  $;HZl��� ������ �2� D�[�h�z������� ԏ���
��3�@�R� d�{�������ßП� ����*�<�S�`�r� ��������̯��� �+�8�J�\�s����� ����ȿڿ���"� 4�K�X�j�|ϓϠϲ� �o�fYo�a�o�o�+� =�O�a�s߅ߗߩ߻� ��������'�9�K� ]�o��������� �����#�5�G�Y�k� }��������������� 1CUgy� ������	 -?Qcu��� ����//)/;/ M/_/q/�/�/�/�/�/��/�XNOCODE� H]e��GkPRE_CH�K J]k� A �� �< ��� ]ee?w?]e 	 <Y?�?�?�Ù?�? �?�?O+OOOaOsO MO�O�O�O�O�O�O�O _'__K_]_7_�_�_ �?{_�_�_u_�_o�_ oGo!o3o}o�oio�o �o�o�o�o�o�o1C gyS���_�_ ����-���c� u�O���������ᏻ� ͏�)��M�_�9�k� ��o���˟ݟ���� ���I�[�5����k� ��ǯ��������3� E��i�{�U�g���ÿ �����ӿ�/�%�� e�w�ϛϭχϹ��� �����+��O�a�;� mߗ�q߃����߹�� ���!�K�A�Sρ�� -����������� 5�G�!�S�}�W�i��� ����������1 gyS��i� ���-Qc =O������ //�/M/_/9/�/ �/o/�/�/��/?? �/7?I?#?U??Y?k? �?�?�?�?�?�?	O3O OOiO{OUO�O�O�O �O�O�/�/_/_�O;_ e_?_Q_�_�_�_�_�_ �_�_o�_oOoao;o �o�oqo�o�o�o�o �o9K_3�� m������� 5�G�!�k�}�W����� �������Տ�1�� U�g�]O�����I�ӟ 埿������Q�c� =�����s���ϯ���� ���;�M�'�Y��� y�����˿e�׿�ۿ �7�I�#�m��Yϋ� �Ϗϡ�������!�3� �?�i�C�Uߟ߱ߋ� ���ߡ����/�	�S� e�?���u������ ������=�O�)�;� ����q��������� ����9K��o�[ �������# 5AkEW�� �����/' U/g//s/�/w/�/�/ �/�/	??�/'?Q?+? =?�?�?s?�?�?�?�? O�?�?;OMO'OqO�O =/kO�O�O�O�O_�O %_7__#_m__Y_�_ �_�_�_�_�_�_!o3o oWoioCo�o�o�O�o �o�o�o�o)S -?��u��� ����=�O�)�s� ��_������o�o�� ���9��%�o���[� ������ß�ǟٟ#� 5��Y�k�E�w���{� ��ׯ�ï��ُ� U�g�A�����w���ӿ ����	����?�Q�+� uχ�a�sϽ��ϩ��� ���)�;�1�#�q߃� ߧ߹ߓ��������� %�7��[�m�G�y�� }���������!��� -�W�M�_ߍ���9��� ��������AS -_�cu��� ��=)s �_��u���/ �'/9//]/o/I/[/ �/�/�/�/�/�/?#? �/?Y?k?E?�?�?{? �?�?��?OO�?CO UO/OaO�OeOwO�O�O �O�O	_�O_?__+_ u_�_a_�_�_�_�_�_ �?�?)o;o�_GoqoKo ]o�o�o�o�o�o�o�o %�o[mG���}�����!�����$DCS_S_GN KeM���w@5a1�0-JUN-22 11:54 ��V�L-18 22�:49g�����? R�:1�����������R�S]����Zo��5�����  9�VERS�ION E��V4.2.10�ϋEFLOGIC� 1Le?�  	����`)�`8��PRO�G_ENB  ⢄ ���Y�ULSOE  >�q��_ACCLIM����s����W?RSTJNT��M�;�5�EMOb����u�
�ݐINIT �M�jזOPT_SL ?	f��
 	R5�75��C�74H�6JI�7I�5��s�1m��2I�*����&�TO�  2�����V.��DEX��dM����-�PATH �AE�A	\MAINPRG\�Y�k��׃HCP_CLN�TID ?� �� *�����؂I�AG_GRP 2�Re ����`E��  F?h F�x E?`��D�y����B�  �Ģ����A�/�Cf�  Cyj�Y�d�Cj�q�B��i���mp3�m6 7890123456���`��  A�f�fA�=qA� � AхA��WHAľ��������A����̱���@���g�ApX�����A���vg�B4�� ���2���
���(�A��A�
=A��B���A��
A�Q�A��������j������j!�	n5��{+A�Z�̶��ZѾ�}������A���������h�zߌ���߰�6�EG�A@���:�RA5Z�/���)��#F�Z� b�������*�<�6؟Pz�AJ��Y�?���9p�A3\)�A,��A&����~������4�}cF�]��AW��UP��J��C��<Z�u4��-Z�%G�� �0�B�T�6�%�
	n ��?Q��%o�w ��Yk�) M_�kc��Q����i�����=�
�==�G��>��Ĝ��7'Ŭ��6�7���@wʏ\&�p�$%���@�Ah��/ A���<i��<x�n;=R�=s���=x<�=�{~Z�;��|%�<'�'�����?�+ƨC�  <w(�U�� 4"w����&����%��\က?ň?� ?6?H?h�$T?~??��?�?�?�?�?�?)�7L?S�FB$��/Eͽ�4OG�ΐ
Ա��iD�5L�x�CA��GX�@j�|�챤��O�L����Oʹ�%_sNED � E�  Eh� DQPXR:_���_����u;Z¨?��s;�a����|;[���
�޳�0y���%ŨP�D�t���O�oC3[H ������s_�_o_o�I�4o:b���Y����u����B����	o�ouo�o�o�o��o�o�o@p�M�?��������h�>���@�2d�=<��=�Du;ě�Pu���CT_CONFI/G S׷񓄄�eg?�ʱSTBF_TTS���
q��s�������v�9�MAU��f�x�M_SW_CFtpT׻�  	�ЊOCVI�EW�pU������Y�k�}������� �rG�܏� ��$�6� ŏZ�l�~�������C� ؟���� �2�D�ӟ h�z�������¯Q�� ��
��.�@�ϯd�v� ��������п_���� �*�<�N�ݿrτϖϰ�Ϻ���\|RC �V�5�r!h���9�(��]�L߁�pߥ��tSB�L_FAULT �W�����GPM�SK�w��hpTBRF �X��>��q�o��F�X���TDIAR	�Yxy��sM!�UD1: �67890123�45��rM!�wh�P (�����	��-�?�Q� c�u�������������@���F��	�"
��<Mt�RECP���
�������� �*<N`r ��������);8/�UMP_?OPTION�p�ޢR!T�s��s%P�ME�uf/Y_TE�MP  È�g3BȈp� �A� �$UNI�p�u�!���YN_BRK �Z2��EDITO�RX!^!�/2_j E_NT 1[��&��,&PNS00�01 OMING� LEFT T_�f2@,&MAI�N ]?o?&PICK_INC�?�@,5&HOME��?�? )&PL�ACE_JACK�PO�4�?�qa&�C@STIC_P�ALLEO�q�&y4OF@RIGH�=��&GRIPP}E�LOSE nO�@&&�EOPE8^ �O@&&K�C�HO�p_&CAL�IBRA[!CHE�CK�0GO�r&C�LAV �C AO@'�&
<S�B�O-[	M?ID_POI@0jO�@*&CAME�A_X E��-[�:LHE�Q_S@*�&MOVETO�1T1t_y&FIND_TOT8F	 N_�r<�0	I�QUo3Ui3 Qb@-o�p�0MGDI_ST�A�%<q�!�q 0N�C�c1\� �P�9~
9~d(/ o������� ��#�5�G�Y�k�}� ������ŏ׏鏀% � �$�6�D�\qD�j�|� ������ğ֟���� �0�B�T�f�x����� ����үL�����'� 9�S�]�o��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� �����1�K�U�g� yߋߝ߯��������� 	��-�?�Q�c�u�� ������������ )�C�9�_�q������� ��������%7 I[m���� �����!�M�W i{������ �////A/S/e/w/ �/�/�/�/���/? ?+?EO?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O�/�O�O_#_=?G_ Y_k_}_�_�_�_�_�_ �_�_oo1oCoUogo yo�o�o�o�o�O�o�o 	5_'Qcu� �������� )�;�M�_�q������� ���oŏ���-? I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ˏݏ� ����7�A�S�e�w� ��������ѿ���� �+�=�O�a�sυϗ� ��#�կ������/� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}�������� �����'�1�C�U�g� y��������������� 	-?Qcu� ������� ;M_q��� ����//%/7/ I/[/m//�/�/�� �/�/�/�/)3?E?W? i?{?�?�?�?�?�?�? �?OO/OAOSOeOwO �O�O�/�/�O�O�O_ !?+_=_O_a_s_�_�_ �_�_�_�_�_oo'o 9oKo]ooo�o�o�o�O �o�o�o�o_#5G Yk}����� ����1�C�U�g� y������o��ӏ��� �-�?�Q�c�u��� ������ϟ���� )�;�M�_�q������� ��˯ݯ�	��%�7� I�[�m��������ǿ ٿ����!�3�E�W� i�{ύϧ��������� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s���� �ϻ���������'� 9�K�]�o��������� ��������#5G Yk}����� ��1CUg y������� 	//-/?/Q/c/u/�/ ��/�/�/�/��/? )?;?M?_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�/�/�O�O �O�O?_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �O�O�o�o�o�o�O +=Oas�� �������'� 9�K�]�o����o���� ɏۏ�o���#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ�߯ 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qϋ�}ϧ� ���������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�ϕϟ�������� ����/�A�S�e�w� �������������� +=Oa��� ������' 9K]o���� ����/#/5/G/ Y/k/��/�/�/�/� �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcO}/kO �O�O�O�/�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o�Io[ouO �$EN�ETMODE 1�]�E� W �@�@�a��D�o�`|hRROR�_PROG %j%F�oy�eTA�BLE  �k��OCUguw�bSE�V_NUM �b?  ��a�p��a_AUTO_ENB  �e�c�dw_NO�q ^�k��a�r  *�*�p��p��p��p�p�+�p��,��tFLsTR��vHIS�s��A�`�{_ALM �1_�k ��D�|@+-�ȏڏ쏐���"�1�_�r�p  �k�q�bg��`�TCP_VER �!�j!�o2�$E�XTLOG_RE�Qh��y��SI�Z��STKߙ��u���TOL � �ADzp��{A ��_BWDG�`�L�H��b1�DI6�w `�EL�x�d�AM�STEP^��p��`��OP_DO���aFACTOR_Y_TUNh�dɩ�DR_GRP 19a�iR�d 	b� ���`��������glrw��qŖ�?�J ���T���f�w��C_�mC���fC@�BB�OY*B���C�U�|�A��\�A�ʪA�UW�@!�@�"��A�^�����w�z����B	���B#e�A����A��]A��ߩB��|�������Ϫ��ұ��*��Y�4!����~�<7`�>�E<�~Ǐ�
 G�0ռ���BB�ԏϟ��pc������߂�`}dC��N<��B�{D�|�@UUT`�UT ߉�$߿ E�� �߀�'�OHcEP]���O��#M�����KA��|�?��� ��:6:�N�,�9-��4�x�
� ��� m-���!�~��T�e���
{FEATUROE b�EH��a�Handl�ingTool ���BEngl�ish Dict�ionary��4�D St��ard����Analog� I/O����gle Shift���uto Soft�ware Upd�ate�mati�c Backup���E�ground� Edit���C_amera��F���CnrRndIm�J��ommon �calib UI�|��nc��Monoitor��tr��?Reliab���DHCP����at�a Acquis�����iagnos�A���ocume�nt Viewe�����ual Ch�eck Safe�ty���hanc�ed����s` F�rt��xt. D7IO ��fiD�wend� Err��QLC��s�	r����  7���FCTN_ Menuy v��*TP Inf�ac@��GigE�Rd\�p Mas_k Exc� g��HTPProxy� Sva�igh�-Spe� Ski���< � mmun�ic@�ons�u�r7	��Sconnect 2	(�ncrRstruH��*0 eWq JC���KAREL C�md. L�ua��g#Run-Tiθ Env](el� +D�sB�S/W���License�s`� Book(System)��MACROs,�?/Offse��%aH� *�� MR�����BMechSt�op�t  (�%i�	�\6x� ��B�>�od�witchȊ?037.6�;Op�tm�?03�fil�`/7g��%ult�i-T�f��PC�M fun:'8Io�%t1DXMRegi�� r�;FriY F�HK�F��Num S�elT5�I�  Ad�ju��N�A	��Mt�atu�A�O[
��R�DM Robot>��scove��8U�ea)@� Freq� Anly�Re�mR0�n��8UDRS�ervo� �0��S�NPX b�"�SNPCliX�^
�Libr���_�� �c4�P�Vo� t7sGsag1E��{� �1��{�/IQ4eM�ILIB]o7bP OFirm(�GnP7�Acc]�e�TPT9X5deln0zo�8a�� 5Hmorqu>�imula��z��fu�0Pa�!Gn\�t��3&�ev.4e� �riq �oUSB port ���iP� aY �vR �EVNTw�pnexcept� yPfDX�u��VC��r��X8V$ ��o��[��S�PSC�eH�S�GE]�S�UI��Web PlV���Q������WZD?T Appl���x�v���GridHQplay�D`I�&�R�r.��`�7�;R�-2000iC/�125L��2D �Gui�pZ����G?raphic�����DV- Path Ctr������v��dv�DCS<p�ckw!��larm Cause/wP�ed��Ascii<��BLoad` \��Uplr��toS���%prityAv/oidM��l����Gu�氯¢8���s2��t����yc��"��@rp~ ��5�os./�cu �z��%�	trans.b�etw.CRLmaOin N��Q.��therNetZa0z���`��ca ��,RA<p� ��(&,0~Q/C�@o�'����L�<�o�89���NR�T���On��e Hel��<E�@�AQ�{tr�ROS ��7�e퇟� ����sup�rt���v�HapA�[����P9k��GiG� t��Im�0F�0X�P��nsp !+�|�64MB DRAMd���FRO�����l�gell���sh��D���c�;��%�p>v�ty�s�B��� r�B��_R�0��� ~�3���hxP���MAIL⋞}�r ��[�CP�R��q�T�1��[��!Adp	.G�X�s����/4Lz�arHQq�Z2�%Ro��+ax��ߏOPT Pؿ�Ac�'`��TX!qpXpSyn.(RSS)TVquir<`��DR��UT��^� (�uesBs�S���]�V�RS6��duXp�[?��Pmi��3DLb�^��w!e��K�`l B�ui)@n�APL�CKV�Հ�CG�UxCRG���D�D@��LS���B�U���K�! /V�T	AT*&B��C*^�X/TCBm/&4/~'x�~'F�/&p~'�
7�u?TEH1?C6�BB7Vi?C6\�
6FP/�7l/
6G�/�7�?�7d?
6H,O
6IAIO�[FHO
6LN�O+%M@O�G�/�G/
6N�OB
6PdOW�?
6R�?B
6SD_rW`_
6W�_8�W_
4VGF�_�UP2��W�O�W�_�VIB@o�VD\o�VF�/��VO�TUT<b0�1�o�f2�o�bTB�GG$b�lr~��� sUI�`|�HMI"r��pon��`�Q�f�or s�>s�KA�RELK��al�TP�Y�c|� SWIM�ESTTr7458918{��|��� ����+�"�4�F� X���|�������ď� ���'��0�B�T��� x������������� #��,�>�P�}�t��� ����������� (�:�L�y�p������� ���ܿ���$�6� H�u�l�~ϫϢϴ��� ������ �2�D�q� h�zߧߞ߰������� �
��.�@�m�d�v� ������������ �*�<�i�`�r����� ��������& 8e\n���� ���"4a Xj������ /�//0/]/T/f/ �/�/�/�/�/�/�/�/ ??,?Y?P?b?�?�? �?�?�?�?�?�?OO (OUOLO^O�O�O�O�O �O�O�O�O __$_Q_ H_Z_�_~_�_�_�_�_ �_�_�_o oMoDoVo �ozo�o�o�o�o�o�o �o
I@Rv �������� �E�<�N�{�r����� �����ޏ����A� 8�J�w�n��������� �ڟ����=�4�F� s�j�|�������߯֯ ����9�0�B�o�f� x�������ۿҿ��� �5�,�>�k�b�tϡ� �Ϫ����������1� (�:�g�^�pߝߔߦ� �������� �-�$�6� c�Z�l�������� ������)� �2�_�V� h��������������� ��%.[Rd� �������! *WN`��� �����//&/ S/J/\/�/�/�/�/�/ �/�/�/??"?O?F? X?�?|?�?�?�?�?�? �?OOOKOBOTO�O xO�O�O�O�O�O�O_ __G_>_P_}_t_�_ �_�_�_�_�_ooo�Co:oLoyoob  H552ocv�a21�eR78�h{50�eJ614�e�ATUP�f545z�h6�eVCAM�ewCRI�gUIF�g�28�fNRE�f5�2�fR63�gSC�H�eDOCVOvC�SU�f869�g0^�fEIOC+w4�f�R69�fESET��g�gJ7�gR68ަfMASK�ePR�XYx7�fOCOB�x3�h�f�p�h3�v[J6�h53rvH$��LCH�vOPLGz�g0�MHCR�v]Sm�MCS�h0�w{55�fMDSW��v�OP�MPR�t?p2�0�fPCMv�R0���p�fw�2�5�1�g51.�0�fP�RS�w69�vFR�D�fFREQ�fM�CN�f93�fSN�BA7w%�SHLB���M��?p��2�fH{TC�fTMIL�h�rvTPA�vTPT�X�EL��w�rw8��g�`�fJ95vT�UT�95�vUE�V�vUEC�vUF]R�fVCC��O��wVIP��CSC��CSG*vdpI�eW�EB�fHTT�fR�65x@�CG��IG�ݧIPGS�RCv��DG�H72�w�9Q�R76�fR8ة�w�b�85rvR6�6b��wR,�R51��w53"�68n�6U6�2�6.�6v7J74�g75b��د`b�<�R5Y�J5�9.�58.�85�5u4��6m�NVD�vcR6y����87j�a4v�p:�i�R7w��pvD0m�F�R;TS��CLI��g�CMS�v?��fSTuY��6��CTO�f�cp�w7qxNN
�NN�vORS���pF�u3��5�HPM�pz�\�?p�fOPI2�t3�ڸ7rvCPR���L��S��7�vSV�SNvSLM�vV3�D��wPBV�A�PL�vAPV�C�CG�fCCRn�C�D��CDL2�CS�BfvCSKCT��CTBަ�T�C�����CҧTC�v��TC��TC��vCTENvs��T�EZvs�ƧTF
�FJ�G��G��^�H^��I�T�CT)�CCTM��� ��N^��P��P��R
�A�T�S
�Wr	2�VGF6�P2��P2��� ��B�D�FvV��VT�g� �fVT�B��VewIH�V�;�K��V��Gene�dvh]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{���� �����/�A�S� e�w���������я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q���  H5�5y�����R7�8��50��J61�4��ATUJ��5�45��6��VCAܢ��CRI�UI����28�NREv��52�R63���SCH��DOCVr��C��869��0��EIO2e�4��R69�ESE�T���J7�R6�8��MASK��P�RXY?�7��OC�O3��� ��3�n
J6��53��H�LCHN
OPL�G��0�
MHCR�O
SMCS��0�55��MDSW�o}OP}MPR�~
{�0��PCM>�R0� ���[51��51,0��PRS69n
F{RD.�FREQ��MCN��93��S�NBAo��SHLEB�*M�+{�^2���HTC��TMILܯ��TPA��TPTX:EL�*��q8���~�J95N��TUT~95n
U�EV
UECN
U�FR.�VCC�<O�.VIP:CSCNN:CSG^���I��wWEB��HTT��R6m�|<CGmKI�GMKIPGS�JR�C:DG}H72���9=+R76��R�8]P�K85��R�66�L��R,R5m1��53�68[�66�2�6,6nN�J74��75�L�����K�R5�;J[59k58k8m<�54n[6[NVD�
R6[P�87�^l4N�; l]+R7XM�; N�D0[F,|wRTS�*CLI����CMS��{p��S�TY;6mCTOh�����7��NN�[;NNn
ORS.; �.l3�k5�[HPM�L,{���OPI�Jkp�\7��CPR�~+L�;S�7n
S�VS��SLM
Vs3DL=�PBVN:wAPL��APV~
wCCG��CCR�CD�;CDL�JC�SB��CSK~CT=;CTBNJېK�TC�*��ΜC>KT�C>���^�TC��TC
CTE��k�n�cTE��k�.KTFޜ�F�GΜG��N�HjN�IN{T��CT];�CTM�M�;���N*N�P�PΜRޜ}|�TSޜW���JVGmF޻P2�;P2�*T���B�D�F>��V��VT��k���VkTB~�V��IH;�V�@��KKVmKGene��~����� +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ��1CUgy �������	 -?Qcu�� �����//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������߀��/�A�S�e�w����STD��LANG���� ���������"�4�F� X�j�|����������� ����0BTf x������� ,>Pbt� ������// (/:/L/^/p/�/�/�/ �/�/�/�/ ??$?6?�H4RBT��OPTN_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�ODPN��	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7I[ m������ ��!�3�E�W�i�{� ������ÏՏ����x�/�A�ted �� z�e�w���������џ �����+�=�O�a� s���������ͯ߯� ��'�9�K�]�o��� ������ɿۿ���� #�5�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߯��� ������	��-�?�Q� c�u��������� ����)�;�M�_�q� �������������� %7I[m� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?�?�?�?�?�?�? OO'O9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �_�_�_�_�_oo1opCoUogoyj99{e��$FEAT_A�DD ?	�����a�`  	zh�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������# 5GYk}��� ����//1/C/�U/g/y/�/�/�dDE�MO b�i   zh�-�/�/ ??"?O?F?X?�?|? �?�?�?�?�?�?OO OKOBOTO�OxO�O�O �O�O�O�O___G_ >_P_}_t_�_�_�_�_ �_�_oooCo:oLo yopo�o�o�o�o�o�o 	 ?6Hul ~������� �;�2�D�q�h�z��� ��ˏԏ���
�7� .�@�m�d�v�����ǟ ��П�����3�*�<� i�`�r�����ï��̯ ����/�&�8�e�\� n���������ȿ��� ��+�"�4�a�X�jτ� �ϻϲ���������'� �0�]�T�f߀ߊ߷� ����������#��,� Y�P�b�|����� ��������(�U�L� ^�x������������� ��$QHZt ~������  MDVpz� �����/
// I/@/R/l/v/�/�/�/ �/�/�/???E?<? N?h?r?�?�?�?�?�? �?OOOAO8OJOdO nO�O�O�O�O�O�O_ �O_=_4_F_`_j_�_ �_�_�_�_�_o�_o 9o0oBo\ofo�o�o�o �o�o�o�o�o5, >Xb����� ����1�(�:�T� ^�����������ʏ�� � �-�$�6�P�Z��� ~�������Ɵ���� )� �2�L�V���z��� ����¯����%�� .�H�R��v������� ������!��*�D� N�{�rτϱϨϺ��� ������&�@�J�w� n߀߭ߤ߶������� ��"�<�F�s�j�|� ������������ �8�B�o�f�x����� ��������4 >kbt���� ��0:g ^p������ 	/ //,/6/c/Z/l/ �/�/�/�/�/�/?�/ ?(?2?_?V?h?�?�? �?�?�?�?O�?
O$O .O[OROdO�O�O�O�O �O�O�O�O_ _*_W_ N_`_�_�_�_�_�_�_ �_�_oo&oSoJo\o �o�o�o�o�o�o�o�o �o"OFX�| �������� �K�B�T���x����� ����������G� >�P�}�t��������� ������C�:�L� y�p����������ܯ ���?�6�H�u�l� ~��������ؿ�� �;�2�D�q�h�zϧ� �ϰ������� �
�7� .�@�m�d�vߣߚ߬� ���������3�*�<� i�`�r�������� �����/�&�8�e�\� n��������������� ��+"4aXj� �������' 0]Tf��� �����#//,/ Y/P/b/�/�/�/�/�/ �/�/�/??(?U?L? ^?�?�?�?�?�?�?�? �?OO$OQOHOZO�O ~O�O�O�O�O�O�O_ _ _M_D_V_�_z_�_ �_�_�_�_�_o
oo Io@oRoovo�o�o�o �o�o�oE< N{r����� ����A�8�J�w� n���������Џڏ� ���=�4�F�s�j�|� ������̟֟���� 9�0�B�o�f�x�����>ȭ  ��ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ �������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/�/�/�/�)  �(�!�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |������� ��0�B�T�f�x��� ������ҏ����� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� \�n������������� ����"4FXj |������� 0BTfx� ������// ,/>/P/b/t/�/�/�/�/�!� �(�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFoXo jo|o�o�o�o�o�o�o �o0BTfx �������� �,�>�P�b�t����� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�D�V�h� z�������¿Կ��� 
��.�@�R�d�vψ� �ϬϾ��������� *�<�N�`�r߄ߖߨ� ����������&�8� J�\�n������� �������"�4�F�X� j�|������������� ��0BTfx ������� ,>Pbt�� �����//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? �?�?O O2ODOVOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����������Ω�$FEA�T_DEMOIN�  Ӥ�����Ԡ�INDEX�����ILE�COMP cw���4����*�SETUP2� d4�>���  N i�'�_�AP2BCK 1�e4�  �)�Ϩ����%��пԠ 7�����ѥ��'϶�K� ڿXρ�ϥ�4����� j��ώ�#�5���Y��� }ߏ�߳�B���f��� ��1���U�g��ߋ� ����P���t�	�� ��?���c���p���(� ��L���������; M��q ��6� Z�~�%�I� m�2��h ��!/3/�W/�{/ 
/�/�/@/�/d/�/? �//?�/S?e?�/�?? �?�?N?�?r?O�?O =O�?aO�?�O�O&O�O JO�O�O�O_�O9_K_ �Oo_�O�_"_�_�_C��w�P{� 2���*.VR�_o�P*oCo�SIomoWU`�PCuo�o�PFR6:�o�nYo�o}kT�$�eN|��x�otVV*.FoD��Q	�c��|a��{STM�+��b��`�V��z��{H G���<���X�j����zGIF	�3�>��܏8��zJPG�����>���`�r��~jJS��:��P͓(��%�
JavaScrgiptf���CSW��=���h� %C�ascading� Style S�heets�\P
�ARGNAME.SDT�|\A�\-���M�]�n��]�DISP*d�G�A����񿀵�򿞿
TP�EINS.XML�!�Ϳ:\5��U�C�ustom To�olbarvϥ�PASSWORD�~z^FRS:\���x� %Pass�word Con�fig�Ϧ���� Y�@���ϥ�W_��{_ ���߱_#��G�Y��� }����B���f��� ����1���U���y��� ���>�����t�	�� -?��c���� �L�p�; �_q �$�� Z�~/�/I/� m/��/�/2/�/V/�/ �/�/!?�/E?W?�/{? 
?�?.?�?�?d?�?�? O/O�?SO�?wO�OO �O<O�O�OrO_�O+_ �O$_a_�O�__�_�_ J_�_n_oo�_9o�_ ]ooo�_�o"o�oFo�o �o|o�o5G�ok �o��0�T�� ���C��<�y�� ��,���ӏb������ -���Q���u������ :�ϟ^�ȟ���)��� M�_�������H� ݯl�����7�Ư[� �T��� ���D�ٿ� z�Ϟ�3�E�Կi��� �ϟ�.���R���v��� ߬�A���e�w�ߛ� *߿���`��߄��+� ��O���s��l��8� ��\������'���K��]��������� ��$FILE_DG�BCK 1e�������� < �)
S�UMMARY.DyG��e�MD:���-q�Diag� Summary�.;�
CONSLOG#q�@�Console� log�:�	T�PACCN�%��1<TP A�ccountin��;�FR6:I�PKDMP.ZI	Pei�
}�=M�Exceptio�n�;�*.DT��/q�FR:\��>.�FR DT Files>/�j MEMCHECCK'��/��Memory D�ata�/��(i{\)�!RIPE�p�/�/A?�#%1� Packet 9L��%�b"1STAT;?"?4?�?� %]2St�atu_/y<	FTAP?!O�?%O�'��mment TB�DNO�'��)ETHERNE�?�&O�!�O�O@Et�hernf0� fi�gura�A�8ADCSVRFBO(O:O�S_�3P verify allV_��$���UDIF�FK_1_C_�_W3mXd�iff�_�W�!PCHG01�_�_�_]o��1�_�o�R�i2 So:oLo�o�_�o�o"b�3�o�o�oe ��o�vVTRNDIAG.LS��BT��!�q O�pe�Ch1 Eno�stic�'�<�)VDEV�rD�A0/��m��1V�is�Devic9e� �IMG�r��H�Z��V3��Imsag���UP6��ES5�ʏFRS�:\5�@/B Upd�ates Lis�tv�;�݀FLEXEVEN�OΏ������1�� UIF� EviAi?�#����)
PSRBW�LD.CM%�e��a�=�x�� PS_R?OBOWELoO9��AIOׯ����'��BNet/IP�pa"��#ߌ)��GRAPHICS4D������%4D Gr?aphicsZ/�'w�' 2GIG?��o���&GigqE���#���2�SMOc����'~P�/Email$��=��\��SHAD�OW��h�z���#�Shadow C�hang���& �~��RCMERR�����ϓ��#X�CFG Error���t��6� �+���3CMSGLIB ��r߄������2��x�����*�)��ZDT�s����'�ZD0�ad9���&=쿢NOTI_v������%Noti�fic�B���&�A�)��u�X�d������������������� ��AS��w� *<�`��+ �O�H��8 ��n/�'/�� ]/��/�/"/�/F/�/ j/�/?�/5?�/Y?k? �/�??�?B?T?�?x? OO�?CO�?gO�?`O �O,O�OPO�O�O�O_ �O?_�O�Ou__�_�_ :_�_^_�_�_�_)o�_ Mo�_qo�oo�o6o�o Zolo�o%7�o[ �ox�D�h ���3��W��� �����ÏR��v�� ���A�Џe�􏉟�� *���N��r������ =�O�ޟs����&��� ͯ\�񯀯�'���K� گo������4�ɿۿ j�����#ϲ��Y�� }�ϡϳ�B���f��� �Ϝ�1���U�g��ϋ� ߯�>ߨ���t�	�� -�?���c��߇��(����x��$FILE�_FRSPRT � ����������MDONLY 1e���|� 
 �)�MD:_VDA�EXTP.ZZZ���z�Q�`�6%�NO Back? file +�B��U�W��A��� ����Q�0��Tf �����O�s �>�b�o �'�K���/ �:/L/�p/��/�/ 5/�/Y/�/}/�/$?�/ H?�/l?~??�?1?�?��?g?�?�? O2O��VISBCK	����*.VD3O}O�0�FR:\L@ION\DATA\hO��2�0Vision VD~�O�8?*.CAM�O_� %	�A�C�O�L�GigE Cam�era Definit�@-_�?}_�? �_O�_�_f_�_�_o 1o�_Uo�_yo�oo�o >o�o�oto	�o-�o &c�o���L �p���;��_� q� ���$���H���� ~����$�I�؏m�7N�LUI_CONF�IG f��|_A|� $ Z��{��ӟ���	��-�;���|xc�e�w� ��������S���� �(���9�^�p����� ��=�ʿܿ� ��$� ��H�Z�l�~ϐϢ�9� ��������� ߷�D� V�h�zߌߞ�5����� ����
���@�R�d� v���1�������� ����<�N�`�r��� ������������� &8J\n�� ������"4 FXj|��� ����/0/B/T/ f/x//�/�/�/�/�/ �/�/?,?>?P?b?t? ?�?�?�?�?�?w?�? O(O:OLO^O�?�O�O �O�O�O�OsO __$_ 6_H_Z_�O~_�_�_�_ �_�_o_�_o o2oDo Vo�_zo�o�o�o�o�o ko�o
.@R�o v�����g� ��*�<��M�r��� ������Q�ޏ���� &�8�Ϗ\�n������� ��M�ڟ����"�4� ˟X�j�|�������I� ֯�����0�ǯT��f�x�������?�x�Robot S�peed 100%������ �2�?��H�x8�E��$F�LUI_DATA g���u��?�g�R�ESULT 2h�u��� �T��/wizar�d/guided�/steps/ExpertT����� ����/�A�S�e�w���ߗ��Cont�inue wit�h G��ance ����������,�>�`P�b�t��� I��-G�uŷ�0 a�H�����u����ps��"�4�F�X�j� |��������������� H�!3EWi{ ��������?������+��&��ri�p����ToolN�um/NewFram�߇�������//)/;/��0x0?/g/y/�/�/ �/�/�/�/�/	??-???  <�;?�����dimeUS/DSTB?�?�? �?OO/OAOSOeOwO��O��Enabl v�O�O�O�O__)_@;_M___q_�_�_F��m?�_�_�?�624�?%o7oIo[omoo �o�o�o�o�o�O�O !3EWi{�� �����_�_�_,��_ ozon�0�}� ������ŏ׏������1���EST �Ea��rn Stand��;�t����� ����Ο�����(�,:��� �?�7���{���Ϻ�Region>�ͯ߯����'�9�K�]�o�����America� ��Ϳ߿���'�9�@K�]�oρ�@�R�y��i����ϟ�bEditor��!�3�E�W� i�{ߍߟ߱�������}��ular 
��� (recommen�)��(�:� L�^�p���������G�������#���~��/acces�� t����������������(C,Con�nect to Network7 n������� �"4K������s��!I�_�Introduct�� ���//&/8/J/ \/n/�/C�p�/�/�/ �/�/�/??0?B?T?f?x?�?�r�u�i��?9��/Safet��O O2ODOVOhO zO�O�O�O�O�O�/�O 
__._@_R_d_v_�_ �_�_�_�_�_Q��?�? �?,o�?\�j�oo�o�o �o�o�o�o�o�o# �OGYk}��� ������1��_�oov�8i#EoWf/current8� ͏ߏ���'�9�K��]�o���D01-J�UN-22 07?:18 AM���� П�����*�<�N�`�r������烏e��ǯ5l ����Yea ��/�A�S�e�w����������ѿ@2022ۿ��(�:�L� ^�pςϔϦϸ������ 
����  �෯ߋ��Month��s߅ߗߩ߻߀��������'�B6/�U�g�y���� ��������	��-���F�� �m�3nA���DaO�������� 0BTfx7�1������ '9K]o�@��R�_��ۯ����Hou�/+/=/O/a/�s/�/�/�/�/�/8�7 �/�/?!?3?E?W?i? {?�?�?�?�?�?�R���O3n"�S�inute�?pO�O�O �O�O�O�O�O __$_��18+_R_d_v_ �_�_�_�_�_�_�_oo*o�?S�Oio�=O��AMP���o�o �o�o	-?Qc u4X������� ��"�4�F�X�j�|�
�������aoÏ�1H�o��NetDon^O�#�5�G�Y� k�}�������ş�Z� �����1�C�U�g��y���������ӯ8a�Co����;�&�r�ipperO�oo�lNum/FraX�s �o��������� ɿۿ����#ϒG� Y�k�}Ϗϡϳ����� ������6oHo�d��&�)9�K�ActiveW�*��������߀�!�3�E�W�i�(�0x0{������� �����!�3�E�W�i�{�  =�������|�ߗ�MacroS�
��w��s~�-? Qcu����|� ���);M_ q������������/.K,������Open\�o/�/�/�/ �/�/�/�/�/?�:� G?Y?k?}?�?�?�?�? �?�?�?OO6�H�/�dO֏�Summary&O�O�O�O�O�O _"_4_F_X_j_ٟ�_ �_�_�_�_�_�_oo 0oBoTofoxo��[O��oO�RobotOp|o
.@R dv����}_� ���*�<�N�`�r� ��������̏�o�o�o���f-5/G/oClos[�k�}��������şן�����2 �E�W�i�{������� ïկ�����4OFI���]��n1��BetMethod"� ��ǿٿ����!�3��E�W�i�,7Dir�ect entr�y of EOA?T datasϱ� ����������/�A�S�e�v��]�RB��U����h$���Btr�aightOffsetv�� �2�D� V�h�z������12}�� Tool�� ����/�A�S�e�w� ��������~���ߤ߄�m%�ߚA��AX ��cu��������21298.4993�GY k}��������/-5�C��?���]/1CY /�/�/�/�/�/?#?�5?G?Y?k?�q	-169.1565o? �?�?�?�?�?�?	OO�-O?OQOcO"/4/���)(O/�Os/�/CZrO__/_A_S_e_�w_�_�_�_�_*95?1.8884�_�_ oo&o8oJo\ono�o��o�o�ouO�O�CDm#�ۣO��)�O���Rotation=wW�ocu����������_1?79.868�?C� U�g�y���������ӏ����	��o�oD%3�AV�oY�-?P� ��ɟ۟����#�5��G�Y��-.2586k�������̯ޯ ���&�8�J�\��<-�g���hK���o�����Rn���/� A�S�e�wωϛϭ�l��-29.4700�������"�4�F� X�j�|ߎߠ߲�q�����������J�"ѿ�tp3Zdir/Tp3z�� X�j�|�������� ������_0�B�T�f� x���������������������o�_Ͱ+�%��Measur�ement/Straigh�O�� ���1CU �&������� �	//-/?/Q/c/"�4F�/j|/We��Nums/New�#sj/	??-???�Q?c?u?�?�?�?j0x���?�?OO*O <ONO`OrO�O�O�O�O�p}/�I�/�O�.��/�,Tool�#Use�O`_r_�_�_�_��_�_�_�_om1 o5oGoYoko}o�o�o��o�o�o�o�op
�OQp�OM_!_�,PartF_�� �����)�;�M�_�b2c��������� я�����+�=�O��a� 2y?���(u�'s/Gڰ�#f� ��&�8�J�\�n�����������71.10������)� ;�M�_�q���������<|/�&B�33������)ɟۙPayl?oad1Cm�V� h�zόϞϰ����������
��EOAT� with tot�=�O�a�s߅ߗ߀�߻��������o Ϳ�O)�S���'ϔy� �����������(�8:�L�^��.Ϡѯ ���������������*<N`˿1z  ?��u�3�2C��  2DVhz�h��Ǡ�no(� ��//'/9/K/]/ o/�/�/�/�v4��/��/ns&��	Advanced�/P?b? t?�?�?�?�?�?�?�?OǠ0xw�.O@O ROdOvO�O�O�O�O�O�O�O_���/�/%_�O_mt%?�Mas�s/Center �Q
_�_�_�_�_�_�_�o!o3oEoWoơ-32.3u��o�o�o �o�o�o�o'90K]tڶ�鿛 �o_�^��^��� 1�C�U�g�y�����\onb2toُ����!� 3�E�W�i�{�������p�w �͏�z),��G"0c�R�xX��R�d�v�������ྯЯ���c�1.5ȏ+�=�O�a�s��� ������Ϳ߿�� �?��C���)��RYϦϸ�������� ��$�6�H��-.1999W߂ߔߦ� �������� ��$�6�0H���SžLៗ�Y�k�}ύRZZ���� �0�B�T�f�x����� ��qo������, >Pbt���i�����x.����p �p�|@�Oas�� ��������'/ 9/K/]/o/�/�/�/�/ �/�/�/�/�(��D?*rt�ϣ?�? �?�?�?�?O!O3OEO \�n�{O�O�O�O�O�O �O�O__/_A_S_?�|�6?�_Z?l?~?rt ���_	oo-o?oQoco uo�o�o��Ə�o�o�o );M_q� ��f_ԟ�_����\�TCPVerif�y/&�Method�J�\�n�������ඏȏڏ쏫lDi�rect Entry��,�>�P�b�t� ��������Ο���xA���=��z'��fy>������ί ����(�:�L����298.4992 O�|�������Ŀֿ� ����0�Bϭ�M�C�?�/���S�e� #��?�����"�4�F��X�j�|ߎߠ߻�	-�169.1565 ����������+�=� O�a�s���V�h�&2�)(����Ϲ� #��_@�R�d�v�����������������a95?1.8884��$ 6HZl~������������Dm�����9���#�W �������/�/%/7/I/�`179.868��w/�/�/ �/�/�/�/�/??+?p=?�x�3�V+�?Oa#�PN?�?�? OO1OCOUOgOyO�O��O �-.2586�O�O�O�O __ $_6_H_Z_l_~_�_O?<a?�5��h?�_�?�?#�R�_=oOoao so�o�o�o�o�o�o�o�`�-29.4700�o 2DVhz �������_�_�S���_5��Z�*oofyMean�������ʏ܏�  ��$�6��o*[�G� t���������Ο��� ��(�:���i�'�ĉ��Z)Y�k�}�ax J������/�A�S� e�w���H�Z���ѿ� ����+�=�O�a�sπ�ϗ�V���z����["�����Introductio��3�E� W�i�{ߍߟ߱����� �ߪE����(�:�L� ^�p�����������������9��R��tutojo�g��Overview����������� ����&8��\ n�������`�"4F ���c���]�Sel�ectT1ModeH�� //$/6/ H/Z/l/~/�/O�/�/ �/�/�/? ?2?D?V? h?z?�?��]o�?�?�`(���Enab�leTeachP?endant�?6O HOZOlO~O�O�O�O�O �O�O�/_ _2_D_V_ h_z_�_�_�_�_�_�_ �?�?�?+oI�$�?�/Joinl`g�_�o �o�o�o�o�o�o (:�O^p��� ���� ��$�6�`�_oo{����'Qo>g�ride_moՏ �����/�A�S�e� w���H����џ��� ��+�=�O�a�s������V�h���ܯ��`�H�oldDeadm�anSwitch ��1�C�U�g�y����� ����ӿ忤�	��-� ?�Q�c�uχϙϫϽπ���Ϡ�ίį&��= ����ResetAlarm��~ߐߢ� ����������� �2� �V�h�z������ ������
��.������[����!M߻ą_J1@�������	 -?Qcu�F� �����) ;M_q�B�T�f���Lo��J2-J6�*/</N/`/r/�/ �/�/�/�/�/�?? &?8?J?\?n?�?�?�? �?�?�?���O1Os�#�cgCarȏ yO�O�O�O�O�O�O�O 	__-_�/Q_c_u_�_ �_�_�_�_�_�_oo�)o;o�?OVo�o�& IO��eO�o�o�o '9K]o�@_� ������#�5� G�Y�k�}���No`o���ԏ��o[A�d_X ��!�3�E�W�i�{��� ����ß՟����� /�A�S�e�w������� ��ѯ㯢�����(�����_Y-Z�w��� ������ѿ����� +��O�a�sυϗϩ� ����������'�����
�T�~����_Rotation� ��������'�9�K� ]�o��@ϥ������ �����#�5�G�Y�k� }�<�N�`߂����o��onc�!3EWi {�������� /ASew� �������������(/�� ��[ALa�stScreen �r/�/�/�/�/�/�/ �/??&?�J?\?n? �?�?�?�?�?�?�?�? O"O��/OOyO;+�file/bac�kup�ddevice4O�O�O�O�O_� _2_D_V_h_z_96�Front Pa�nel USB (UD1)�_�_�_ �_�_oo)o;oMo_o\qo�o  EB�CA�OaO�o��%�O�Fi�rectories�o1CUgy@�����>1�P�:\\BKUP_�12-DEC-1�8_01-48-30\\��-�?� Q�c�u���������Ϗ �mJO�o�o$�B��oE�defڏo������� ��ɟ۟����#�:5�Image B �B+�\�n����������ȯگ����"��m��=@'�	�k����A%gripper�P$ToolNum .���ѿ�����+� =�O�a�s�6?�ϩϻ� ��������'�9�K� ]�o߁�DOR�d��������S!G��Typ �O�%�7�I�[�m����������Single �ѝ��� ��*�<�N�`�r��� ���������lg�o���!�g��Comment/cmt�� o��������#����L^ p������� //$/����#�g/-�?���Summary*/�/�/�/�/ ??+?=?O?a?s?�� �?�?�?�?�?�?OO 'O9OKO]OoO��@/R/ȜO�O�!"�/�eprogres_%_ 7_I_[_m__�_�_�_ �_�?�_�_o!o3oEo Woio{o�o�o�o�o�mA�O�O�o�",�O�M�F6�or�����������\-#�I�[�m������ ��Ǐُ����!�8/��of�(:Lss7&�Ɵ؟���� � 2�D�V�h�'�0w��� ����ӯ���	��-� ?�Q�c�u�4�F�X���8|�����ss8z�� ,�>�P�b�tφϘϪ�����\Initioaliz�� B�" ����'�9�K�]�o� �ߓߥ߷��߈�������,	9KIO/s1��a�s���� ����������,�O� D�V�h�z���������@������
�B
�߀�A��]�1�C�2 "�����! 3EWi(���� ����//(/:/ L/^/p//A
O�/��N!��Commentv/??/?A? S?e?w?�?�?�?�?�_ �?�?OO+O=OOOaO@sO�O�O�O�O�M�/���O_�/� �O S_e_w_�_�_�_�_�_ �_�_oo�?=oOoao so�o�o�o�o�o�o�o#g�O�O;e .o������ ��!�3�E�W�i�(o ������ÏՏ����@�/�A�S�e�v�Jp kE����{���� �(�:�L�^�p����� ����w�ܯ� ��$� 6�H�Z�l�~������� s��������͟2�D� V�h�zόϞϰ����� ����
�ɯ.�@�R�d� v߈ߚ߬߾������� ��׿���]�τ� ������������ &�8�J�\�߀����� ����������"4 FXj)�;�M��(�-_�!MacroNumA_ $6 HZl~���s� ���/ /2/D/V/ h/z/�/�/�/�/�O���/?�!��ea�surement �/W?i?{?�?�?�?�? �?�?�?O�/OAOSO eOwO�O�O�O�O�O�O �O_�/�/�/4_^_�� %?71Weight��_�_�_�_�_ o o$o6oHoZoO~o�o �o�o�o�o�o�o  2DVh'_9_K_��y_�W�_��� 0�B�T�f�x������� moҏ�����,�>� P�b�t���������{ ���s�(�:�L�^� p���������ʯܯ�  ���$�6�H�Z�l�~� ������ƿؿ���� }ߟ�S��zόϞ� ����������
��.� @�R��c߈ߚ߬߾� ��������*�<�N� `�ρ�Cϥ�g����� ����&�8�J�\�n� ���������������� "4FXj|� ��q������� 0BTfx��� ����/��,/>/ P/b/t/�/�/�/�/�/ �/�/?�%?�I? ?�?�?�?�?�?�?�?  OO$O6OHOZO/~O �O�O�O�O�O�O�O_  _2_D_V_?w_9?�_ �_qO�_�_�_
oo.o @oRodovo�o�o�okO �o�o�o*<N `r���g_�_�_ ���_&�8�J�\�n� ��������ȏڏ��� �o"�4�F�X�j�|��� ����ğ֟����� �'�Q��x������� ��ү�����,�>� P��t���������ο ����(�:�L�� �/�A���e�������  ��$�6�H�Z�l�~� �ߢ�a����������  �2�D�V�h�z��� ��oρϓ�����.� @�R�d�v��������� ��������*<N `r������ �������G	�n �������� /"/4/F/W/|/�/ �/�/�/�/�/�/?? 0?B?T?u?7�?[ �?�?�?�?OO,O>O PObOtO�O�O�O�?�O �O�O__(_:_L_^_ p_�_�_�_e?�_�?�_ �?o$o6oHoZolo~o �o�o�o�o�o�o�o�O  2DVhz�� ������_��_ =��_�v��������� Џ����*�<�N� r���������̟ޟ ���&�8�J�	�k��-������/wi�zard/gri�pper/ste�ps/SummaryU������/� A�S�e�w�����Z��� ѿ�����+�=�O��a�sυϗϩ�   _�������W���ˡ�TCPVerif կ<�N�`�r߄ߖߨ� �������߯��&�8� J�\�n������� ����������C�]�i"�ˡG IO&� �������������� 0B�fx�� �����,>PW �%�o� _�����//,/ >/P/b/t/�/�/W�/ �/�/�/??(?:?L?�^?p?�?�?W�i�w ��?�O"O4OFOXO jO|O�O�O�O�O�O�O �/__0_B_T_f_x_ �_�_�_�_�_�_�_�? �?�?;o�?boto�o�o �o�o�o�o�o( :�OKp���� ��� ��$�6�H� oi�+o��Oo��Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ��Y���}�߯���� *�<�N�`�r������� ��̿޿𿯟�&�8� J�\�nπϒϤ϶��� ���ϫ��ϯ1���� j�|ߎߠ߲������� ����0�B��f�x� ������������� �,�>���_�!߃��� Y��������( :L^p��S� ��� $6H Zl~�O���s�� ���/ /2/D/V/h/ z/�/�/�/�/�/�/� 
??.?@?R?d?v?�? �?�?�?�?�?��� O9O�`OrO�O�O�O �O�O�O�O__&_8_ �/\_n_�_�_�_�_�_ �_�_�_o"o4o�?O�O)O�oIC�$FM�R2_GRP 1�i�e� ��C4  B]�KP	 KP�o��l�`E�� �o��G[�`OHcEP]���O��#M{��-qKA��}�?pIEl�`:�6:N�uq9-��}u}A�  ��{BH�cC`}�dC��N�qB�{�uEl�d����`@UUT�UT�}�R��a>FD��>�d�>D��=�=��1�U�op�H$:���=:��:.��	:sf�:�Uf1���}�����ۏ����8�KW�b_CFG� j�kT �C�������J�NO ��jF25�3267 973�7K�RM_CHK?TYP  �aKPp�`�`�`�aROM���_MIN��KS���+���pX�`SS�BZ�k�e �fX�KUO�x����P�TP_DEF�_OW  KT|�c��IRCOM������$GENOV_RD_DO �VQnݭTHR � d���d�_ENBϯ ��RAVC�cl�A�L� ��f���`�}EӤ��G
�F�/lG�,�t���KR��`!��vث��r��C�OUZ�`r�l KP�h���e<(�[5��ۿ-�^���w��z̉��h��^�<.�����*���Z���C����,x�Dj>->KQC����W��d����B�`��B��a����i ɑ�D�SMT­csQ��`N����$�HAPTIC_C�NT 2t�e�[�
!���@W�vKSs<x�A�KS���x�C�s2]x�I�KS����H���s^@�x�E�Ԥ����m���>\x�G�������x�<���'�nx�p�KS^X�FEAT  g�Z�� <�8��B�8T�c�X�OST_�\�s1u�iM��V_k 	������2KV��HYe��� $�6�H�HZ �y�����������f�	ano?nymous��(:L ���� �����h��� Z�7I[m��� ������/Vh z��{/��/�/�/ �/�/.??/?A?S? v/���?�?�?�?�? */</N/+Ob?OO�/sO �O�O�O�/�O�O�O_ _8O9_�?]_o_�_�_ �_�?�?O"O$_�_XO 5oGoYoko}o�O�o�o �o�o�ooB_T_1C Ugy�_�_�_��o �,o	��-�?�Q�� u��������Ϗ� ��)�;����� ��̏�˟ݟ��� Z�7�I�[�m����؏ �ǯٯ����V�h� z�����{�����ÿ տ�.���/�A�d� RϬ��ϛϭϿ���!��w�Eb�1v���  P!e�#�����N�=�r�5ߖ�Y� ��}��ߡ������8� ��\���C��g�y� �������"���F�	� �|�?���c������� ����Bf) �M�q��� �,�Pt7I��m����Q�UICC0��!�192.200#.1B &/(1O/+/G!1G!E/V/2�/�{/��/!ROUgTER�/�/!
�$�� ?�PCJO�G???!?!1�68510�/#CAMPRT�?k?=#�111�0�?�6RT?�?��?-O��NAME �! �!ROB�O�?5OS_CFG� 1u � ��Auto-started6�/FTPA��AX� Z��O��_'_9_K_]_ ���_�_�_�_�O�_n_ �_o#o5oGo��O�O �O�o�_�O�o�o�o �_BTfx��o /������� 1�C�U�����o���� Ώ����(�:�L� ^����������ʟܟ �5�G�Y�6�m�Z��� ~�������{�د��� � �C�ů?�h�z��� ������	��-�/�� c�@�R�d�vψ�O��� ��������ϙ�*�<� N�`�r߄�˿ݿ��� ���7��&�8�J�� ���������m� ���"�4�F��ߟ߱� ������������� ��BTfx��� /����a� s���3������ ����/(/:/L/ op//�/�/�/�/�/�pOD@_ERR �wNJ�/�&PDUS_IZ  | ^���4>,5WRD� ?�E^� � guest|&l?~?�?�?�?�?�=DSCDMNGR�P 2x�E0�^| wd|&�KD	P01�.00 8C �  A  %�  

@�?@}�D�9 �������������hg@1g@�����XSM  �?G_�  �P�SO��ygG�E����R���{O��?@�@�D�0
�ZD�O�{g@��@U-w@�k@ew@��O+�+X�I0�+Sy*�d7OIO[OmO�;_GWROU�0y9@��2	�1.C�XQU�PD  Z5��T�PTY�`=�� TTP_AUT�H 1z; <�!iPenda�n�7Hnmai�>kVP !KAREL:*HoQocm�KCxo�l�/mc�VISION SET�P�o�oig�o�o '!nEW�{�����mbdCTRL {=&BD|!�x *�F�FF9E3�\�FRS:DEFA�ULTV�FA�NUC Web �Servery*
�ZdT?f4123456�6΁�ԏ�����}� WR_�CONFIG �|�; oV��!I�DL_CPU_P5Cu�|!B�_��� B�]��MI�N��D1 >zUL~��GNR_IO1�:2| 8��NPT_�SIM_DOΖ�6��NSTAL_oSCRNΖ ��X�INTPMODN�TOL�؛��RT�Y�ݖ�``EN�B��R|�OLN/K 1};h0�����į֯������M�ASTE͐�^��SLAVE ~?�;�RAMCACH�E*�"�OaO_CcFGl�����UO`�n���CMT_OPpu�В:³YCLk����o�_ASG 19�7F1
 �1� C�U�g�yϋϝϯ��π������	����N�UM939
��I�Pi�{�RTRY_CNͿ����Q93����5 ��������J�\0��\0��P_M�EMBERS 2Y��97P $������}��(逐R�CA_ACC 2���[  T�9�`�� 6�)�|"� | |!v��7:�  �b �8%0� !�� ,��|"��X�BUF0�01 2��[= �5 u1u1 � 5 ��@��`uW2u2�������U������6��6 ��6�6`1�u3�uP�6 �6(�6�Z�7��7 Y�7��7P�8 t�t���� �8�8`u�5u5���u6ufӀ8���(�8�Y�9 ��9 �9�9�P�9yd�d� [ 1�1�Y�1(�U10�2��2 �2��2P�2�2��2�(�20�3��3 �3��3`u4u�3��3 �3(�30�4���4 �4�4P�4*�4 �4(�40���2�� ���	�� -�?�Q�c�u������� ��������); M_q�����	��3��HQ2 22!2)21 292
4H��4X ��a��i��:4x�� �HQ��2��2"4� ������"4��� ������B4�HQ� �24��2j4!HQ! B BB4(!HQ0!5B 4@!5Bj4P!5BY 5B B4h!HQp!uB4�!uB � uB24�!uBB4�!HQ �!�B4�!�Bj4�!�B0:4��花2��]�P4�<�HQ��<HP+T�.QВX�HIS���[ �v� 2�022-06-1�2{� ��.Qdt�ЃRka8 ��2��S(�ST�P&�  ?8�T9` �S&��_�_�_oo+o���ʿgY�Pv_��9�r�_�P ( !Ѝ��R�Pga`�P# g :�Pga^@mc;"H� ]��.Q�cX�d`  ' � ChF Z�p�Tx  :�a��b�* ��T���c[�   .W ��T��T��d��md��TT�Bi0U9Pl;3�c��4�ЕV�P�`#t`�a`�P�aYOb.P�P,R�` Kr�`;r��gb�`�R�`H�R�`;qb�h�a^�`Kq"�`�b�`�r�`;r��`!  6�ld0p�Rp�bT�zhr�To�c�P,Rt`7 � \�TS�P  ��R�`�R�`�R���r�x�`*�`�R�`P/��`�R�`>�4�`P;r�`�R�`�`�'JpA�` / �p�Rp % Y'p;rT�z7��Srdh�rt`;r�P/�[`�`6 
T��R�`�3 	 T�`Kq$ �`�b�`�b���m�u+������`5��Xp)R�`Ep�av�zT�2�a��,��Ilh�/���B���xtb����rd�:s�h�r��.���N�`Sr�`/��`	"o �ofc��pCqWT�z�2�gb��U/��O�P��2t`E-1PL�Pǂ�P��	/�PC�U�`�b�`�b8���`��3�hג���c��,R�`1  R���bd��b�`[rt��� uCY� R_d_ 
��p�R�p�P��tb�p �P���P���R�p�R�p .o����,�>�P�>o������`�P;�a��; �aͽL��pT�����r�p�`���`9�a�b�p ���c���b�p���p�` ��d��p�b�pr�p�r �pr�pwϭ����� ����`�t��u��A��� ��	��`�+�=��T� f�xݤߟ��`�Ȥ� �������:��qՏ 0�B�xߊߜ߮ߌ��b ]���������^1ޱ���ѓ ���Wq8�J��d�����4��������7�:ha�����/� S��`���`Q�� u���1�CY� Xw���
�,� Q��� �(�0 3,ݭ3�9`�	/ /-/?/Q/c/u/cϾ���"��"��"�Q���"�� Q@�$�H ,� QP ,�� QX�$` ,�� Qh ,� Qp �,� Qx4�4�^4� ,� Q�/4U����������`�A�������2���p��2���2� �2� �2� �*�$��$�4�
4�2�0�20�2&0�*4� 24�">0�"F0�"N0�" V0�"^0�"���`� aB�aB�aB�aB����B� �B� �B� ��$�B� �B0�B0A�4�B0�B&0�*4�24�B>0�BF0�BN0��BV0�B^0�B����"���ER���UR �UR�UR� UR� UR�� UR� UR� UR0� 
4�R0�R0�R&0�R.0�24�R>0�RF0�R N0aBV0aB^0aB���Af�b�b�l� 1b�1b�1b� 1b� P1b� �`�"q�$s4At
4yb0yb0v"4w*4�b60y:4�bF0T�bN0R4�Z4��"��_��b��b� �b��b��b��b�  �b� �b� �b� �� @�0�0�0c4 er&0er.0er60er>0dB4�rN0bV0b^0�bh�I_CFG �2�� H
�Cycle Ti�me!Bus|�b#Idl�r^�tmin|+��Up�v�qR�ead�wDo�w������sC�ounya	Num �r�s�|+�� yZ�h�PROG�r�����)�/softpar�t/genlin�k?curren�t=menupa�ge,1133, �����/�
�"h��SDT_ISOL�C  ����;��$J23_D?SP_ENB�e�����INC ����#s�A	 ? �=���<#�
r�>͙:�o ؑ�`�!�+��OB���C�������E�G_�GROUP 1��e��< A���͑~)��3�?(��Я Q����/��S�e�w���'��=�G_IN_A�UTOR�����PO�SREM�_�KANJI_MASK��׺KARELMO�N ����"y N�g�yϋϝϯϲ�%�J�������$��|쿢�KCL_Lǰ�NUM���$KE�YLOGGING���UQd����LA�NGUAGE ��m��DEFAULT {�6�qLD�q�����P�F�����G�Ҏ�����3 u�� � '�' + � ; >�L��;��
$�(U�T1:\��D�  F�S�e�w�������������(
FRA:\RSCH2����LN_DISP �����㯹ԟOCTOL��!D�z��n�ɑ��GBOOK ��ݕq����p��	 -?Qcs����	a	���ٍ�H���<�Ñ��_BUF�F 2�e� �2���M�0 �L^����� ��� /-/$/6/H/�Z/�/~/�/�/���DCS ���ёB��	����#;_���
��B�wN��Z2��8�j%>@B�5�A��B��B��5A�ab��� I�O 2��� �p�?�p���?�?�? �?�?�?�?O$O4OFO XOlO|O�O�O�O�O�O��O�O__0_D_��~�ER_ITMb�d���_�_�_�_�_�_ 	oo-o?oQocouo�o �o�o�o�o�o�ok9NtPSEVΰ��nVTYPb��_m8�}�RST$��%�SCRN_FL +2�}=�������)�;�M�_�q��T�P:�b�\r��NG�NAM����m��$U�PS`�GI�p������_LOAD�J�G %��%DF_MOTN���1���MAXUALcRM!�� 瞕9
E��_PR��� ��E�Cc�����k7��k�P �2��� �$	V���ΰ�ΰ#�� B���$��!�Z��H� ��t��������ί� �+�=� �a�L���h� z�����߿ʿ���� 9�$�]�@�Rϓ�~Ϸ� �����������5�� *�k�Vߏ�z߳��ߨ� ��������C�.�g� R����������� ����?�*�c�u�X� �������������� ;M0q\�>��DBGDEF ���������� _L?DXDISAˀ����1E�EMO_AP�ŀE ?��
 ���0BT�fx��E�FRQ_CFG ���m�A ��@����<��d%�/�t�ؒ����*T /V" **:_"��R/d(� ���/�/�/�/�/�/�/ ?5?���^?TPO?�?s<�=�<,(3?�?�� �?O�?+OO<OaOHO �OlO�O�O�O�O�O_�_�O9_;�ISC 31���E  ��?�_ ���_��_�_�_E_�WR_MSTR ��-}eSCD 1���_fo�_�ouo �o�o�o�o�o�o, P;t_��� ������:�%� 7�p�[��������܏ Ǐ����6�!�Z�E� ~�i�������؟ß�� � ��D�/�T�z�e� ����¯���ѯ
��� �@�+�d�O���s��� �����Ϳ��*�ϰN�9�r�oMK��&m���$MLT�ARM��9'�� x3� ����>� METPU� R���.iNDSP?_ADCOL�� ��CMNT1� �$�FNM�Q�"�FS�TLIr�c�` �&n���������$�_POSCF��\��PRPMP���STv/�1�&k 4�#�
a�v1a�q�� ]���������� ����A�#�5�w�Y�k������������$�SI�NG_CHK  }u�$MODA���_[�˯�DE�V 	�
	M�C:QHSIZE��P�TASK� %�
%$12�3456789 ���TRIG ;1�&k l���~9M~=�YP�~53EM_�INF 1�9+�`)AT&F�V0E0R�)��E0V1&A3�&B1&D2&S0&C1S0=�)ATZ�/$�H!/I/�=q/ (A�y/�/\/�/�/�/�/  � ?���	/z?-/ �?�/�?�?�/�?�?O .OORO??�O;?M? _?�O�?�?_=O*_�O �?`__�_k_�_�_mO �_�O�O�O�O8o�O\o �_mo�oE_�oqo�o�o �o�_�_F�_oo ��So��o���o ��B�)�f�x�+�� Oas�����,� c�P��t�/�������|ΟJNITOR���G ?e   	EXEC1iê�2�3�4�5��� �7�8�9i����|��|�"� |�.�|�:�|�F�|�R��|�^�|�j�|�v�|�2���2��2��2��2���2��2˨2ר2��2�3��3��3�"�R_GRP_�SV 1�� �(������k��
�����"��x|��1��_Dm��~׳ION_DB' ��+c�  ������D� "Zc�#)��l��l���DĐN   E��]��)������D-ud1: RSCH\ݟ�ϰ��"�PL_NAME� !����!�R-2000i�C/125L, �Handling?Tool  \�"��RR2�� 1��(�@��R� d��'�9� K�]�o߁ߓߥ߷��� �������#�5�G�Y� k�}���<2#��� ������&�8�J�\�n�<<��������� ����(:L^���|�  �����  �� � ��  A� W B� T� ����
� �� ��� g ��� � B� �z� �  C��C���P E;�� E@ D�����D� ��� ����]���
E��)>g+E(� :9Z�H�%Z!fn/W}� �Y"JJ� =D����>>�+���(#�P0'%��(/2!&!F!b%J!% 2%F%F!&!%f6)�%
J!m� N+2%J!& �!�J2(��$I"�,1&S�)?$?0'0� �� a2��h?n1 b1F%n?�3F!�� f4&!�=�g� �3�1�f?�3�`�3�?�6Fp E"B�?�3�4F�?}6>BO|7��bO�N� E#��E��E��r"����  � �O�K��d�C�D�O Y �O"_0W�@��B]S�ǇW%n__�_KVc �X�_�ZAp� =��S�����_�_T	o�W��P��TB�@i���Wogl���U�	`�_�o�o�o}a:�oA���o�o~;`\�)r�=f�_ O:w|�l~{�_�X��������RN�� 1���R��bl6 Ē��w�@�%?|� v���?��<v���@�6�Z1�z��;�	l��	�  ~�� �,^{�|������ � s? � � �䂱��K�l,K����K��2KI+��KG0�K �U�����O=���@�6@ t�@?�X@I�b�������N�����
��ՙ��G��_�����v�~1a��k�ô� �"���  �X��ￒ4������r���  ������bW|��>�T���f�����	'�� � ��I� �  ��Q��:�ÈƯÈ�=���ޥ*�@����`��*�`��e4��[�p�  �'��S���?��ab���^���C��MB� C4� ��B"tʱ����}�α��� � � �J�����B�P �*u�m&p�F��� k�	���zϳϞϰ����5~ ������� �,0�:�d  }��?�ffA_$�6��� w`k�}�b+�80��ߡ�?�RI�����(0���P�؀���΃΄8������Qa;�x5;���0;�i;�d�u;�t�<!�!��C�R߄�`����&p?fff?�?�&��Nd@��A�#��@�o[ ��0��{���v��� t���d纄U�*��N� 9�r�]�������������0���F.p��, ��P��q��C�?MEtPC�3�1�3� ���<'` K]���`�� ���g-/�T/�x/ �/�/�/M��/�/o/?��/,??P?;?�aA!�x4�P�R�?AJ?�?�F8A�/C<?��`�?�?OO0������W0OC�T��`G Ca-O*�4��0��1�Ab�ܮ���b�C@_;CLn��BA�Q��>V�.È�����Y�\ϼ��
}OOc���Q��hQ�@��G�B=�
?h����O/`���W���ɰ�B�/
=�����Ɗ=2MK�=��J6XLI��H�Y
H}���A�12ML��jLLPB�hH:��HK��n_�P	bL ��2J��H���H+UZBu2O�__�_	o�_ -ooQo<ouo`o�o�o �o�o�o�o�o; &8q\���� �����7�"�[� F��j�������ُď ���!��E�0�U�{� f�����ß���ҟ� ���A�,�e�P���t���������ί��G�ϭ�� C�a|�?;� Ĉ��]��d�CVF酿���xI[Կ�@��Kտؿ� 
E�� �ƿ�K��@(�A�_�h�M����~����N��nπϪ�3lCq��ϬϺ¢�����ϰt�.3���}���k���q?'�3�JJ�ـ^�L߂�pߦߔ��5P>�P�����T�`�7�"�[�F��a�h�����{������  fU���%�� I�4�m����������������
���)Z,  ( 5�{0HB�~����  2 �E�G!�3E�Lݏ��q�5B�X�0w1Q�C�l@�1  @Q�L�0 k�}�b��6��}Ӥ���/L///?�@#�8�4�y�0e��4�;
 0/�/�/�/�/�/ �/�/?#?5?G?Y?k?�}?�J�2����V{�H��$MR_CABLE 2��ؿ ���T&��@P@PA? PA��1�1�  ´� �0C�06!O4>ߔB�l�Y�=� #�2M1?l�� �����?~�6�,  �� �( l6#N�/H�B��:�{m�� �G"M����BZx,O>L<�N@` �L�D���B��CB��  �� B?Ϝ͸�]�E�? �3�O���O��O�O_ _ _�_�_V_�_z_�_ �_�_�_�_�_o
oo@�o|oRo�o�dE���  B��0�B�B�^�B�A(B�,��B��B����B���B��v�B��}B����B�|!B�c=�B�FB�.��B�zB��R�B���B����B����a�}����@���������� ������`�� ���7p�;p�?p�Cp��Gp�Kp�Op�Sp��7p�;prOpx 2026/0��|5*�3OM ��9����K .���%% �2345678901��u ���qR6 �6 ;6 6!�
�w�mno�t sent *�K�6!�W���TESTFECS�ALGR  egD�;d��a!�
��� ��ЭD�3�l���ŏ׏� 9UD�1:\maint�enances.�xmYD,��kp*��DEFAUL�T��2GRP 2���z  p �5�*N6& � �%!1st �cleaning� of cont�. vG�ilat�ion 56��Bԓ�@ޑ��+�a���"�4�F��m��H��@%��me�ch��cal c�heckW�  ����C �������֯����[���o���roller�������ů�����п�1�Bas�ic quarterlyD�W�i��,��V�h�zόϞ�)�cMw���6 "8��!6 �����M�"��4�F�Xߧ�6!%C ;����ϸ���������
��k�}�Gr�ease bal~�r bush+���}���ߪ����h��/�A�C��geu��.L�t�y��  	3d�2� :�A��	��n���������}��
�gG��6&f�B��-6 ���]�@2DVh��}�
��cabl��6"�� ��@���
!� ,>�������������/}�Overh�au�ϕ�@" !x�J!Q/���~/ �/�/�/�/�$o/�/�h�o? m/B?T?f? x?�?�/�?�/?!?�? OO,O>OPO�?tO�? �?�?�O�O�O�O_SO �O:_�O)_�O�_�_�_ �_�__�_ oO_$os_ HoZolo~o�o�_�oo o�o9o 2DV �oz�o�o��o�� �
��k@���v� �������Џ�1�� U�g�<���`�r����� ����̟�-��Q�&� 8�J�\�n������� �������"�4��� X�����˯����Ŀֿ �7����m�ϑ�f� xϊϜϮ�������3� �W�,�>�P�b�t��� ������������� (�:��^�߿ߔ��� �������� �O�$�s� ��Z���~��������� ���9�K� o�DV hz������� 5
.@R�v �������/8/�\	 T/I/ [/m/��/��+�-�/ �/�/�/�/�/<??? V?H?�?x?j?|?�?�? �?�?�?8OOORODO �OtOfOxO�O�O�O�O�\ ̼?� ; @\ z/Q_ c_u_\=_�_�_�_\w*�_** Q V�P�Oo,o>o obo8to�o�o���� �_�o�o�o�o1C U�o�o�o)��� �	��-�w�� u������m�Ϗ�� =�O�a���M�_�q�3�@��������\\��$MR_HIS�T 2�U��� 
 \d$ 2�34567890�1$�,���R#�9 ]����L�~�[ݯ� ���ʯ7�I�[��$� r�����l�ٿ����� ƿ3��W�i� ύ�D� ����z��Ϟ����� A���e�w�.ߛ�Q� ��SKCFMAP � U���R��Q��߳�ONREL  ���������EXC/FENB��
�Ӳ���FNC��JO�GOVLIM��d��g��KEY��zj�s�_PAN�ظ����RUNZ����SFSPDTY�P>�	��SIGN|���T1MOT\�����_CE_G�RP 1�U ���4 �_h�Q�U��� ������x������� ��?��4u,�� b����)� "_��|�p����/��PD�_THRSHD { Q�F@ )�QZ_EDIT�������TCOM_C_FG 1���!�؏/�/�/ 
p!_A�RC_���I�T�_MN_MODE����)�UAP_�CPL�/-�NOCHECK ?��/ �� M?_? q?�?�?�?�?�?�?�?�OO%O7OIO[O��N�O_WAIT_L���e'/�ODRDS�P�#��)�OFFS?ET_CAR[ �/��FDIS�O�CS_�A� ARK��f)O�PEN_FILE��@��!f&� OPT?ION_IO{���QPM_PRG �%��%$�_�_-SWmOP�?���������U����  ���GQ��P'�Q	 �Q��QQ��zD��@RG_DSBL  �����No��ORI�ENTTO��?"Cٴ����A �BUT�_SIM_DYW������@V�@LCOT �����Q��$dQ�Z�dIe�a<Q�`_PEX� �On�dRAT�' d)���d�@UP ��m�!ݐ�QcI���y�$PARA�M28��(��@�c �`/����%�7� I�[�m��������Ǐ ُ����!�3�E�Q�2�t���������Ο �����Q�<c�@� R�d�v���������Я@����������O���  ��  ���  A�  �BC�[ B�{s���3�H7��  �Y�?�>�BC�zC���z`yaQ�P �E;� EE D�	���M�Dn�����n������  �������E���Ѳ�gӳEc(�ȳ��Z��@Z�Ͷ�ɲ��/�� %�2�B��ʱ��b�Ȳ�>̅Ζ{���m�Ӱ���ÎP���ū���������
� ���������������(��2���m��NӰ�� ��ε^т���ȕ�������Bٮ�̳����ǂ�}���	��Ȁ��
����<����Ѓ����:���� 0l�n��l��`��~�>h�Fp Eʰ�����v�F3�%�� ��$炱
�4�+�0�&AB�g�y��d#�����������J�J�-CW%P�@��`X4^T
Ap?��g����q[�� ��BZ��2 ��P�mB3	`�HBTf%:��o�a����3 B�`�Z��2�� �Q/&+(I/ /m//�j/�/�/�/�F�r�pO�7p1�!�(�!���t0l�6!dA`��� @��?>�"1�G�?m@"1xb�˴x�"�P>;�	l22�	�P *0� ��,^�P�Pk0��� � s �� � ��2� H���9H�H���H`�H^yH�R�,�hW��?�<� C`B�C�ʰC4D;0O�#�9W�� ��k��}`�ʰ>A"O4O�FO�#�B<�{��KA��)O �"j��OK@���C�'$/2�?��? Q�V�/�0_�%	'� �� NRI� ��  ��MJ=����r_�[R@��_�P�N"a�_8["b�/�O�'N�`o  !'�`4d�1[@B:�B�}`
BoOAoSo -� O }�
A�8��`%�>�B�&B� �f ����Q�e���/��/;&_J\pOU�5``P�u�a�u E,KB:z�b�1�D�?�ff�����t �)�[q8XK@?�M�?��.1Rz(K@{�P���y�1�z3z4�Sj����Zq;��x5;��0;��i;�du;�t�<!�ڲ?���04�S22�?offf?�P?&,��Wt@��A=#B�@�o[J�KI �b'���[p"5�� 7�� �f4�֟������ 	�B�-�f�x�c����� ��ү����m������4P��E C�۴r���?�����Ŀ��� ӿ���	�B�-�f�/ �ϕ�W�M?���7� � s�$�6�H�Z���o߁߀ߴߟ�����������A�$� �6�C���[���텹���?Ƀ؉�����KI�mرS�W��C� p�` Ca���ʣ����F�@I��Zn��bC@_;�CLn�BA�Q�>V���È����Y��\���
�)�����Q��h�Q�@�G�B=?�
?h�â�� ���W����ɰ�B/
=����Ɗ=JM�K�=�J6X�LI�H�Y
�H}��A�1�JML�jL�LPBhH:���HK�, 	�bL �2J���H��H+?UZBu�� ��|������ !1WB{f� ������// A/,/e/P/�/t/�/�/ �/�/�/?�/+??O? :?L?�?p?�?�?�?�? �?�?O'OOKO6OoO ZO�O~O�O�O�O�O�O _�O5_ _Y_D_i_�_8z_�_�YGϭ�_�_� C�a3��_ �爓�	ooCVF��1o8o����o�P���K�o�o� 
AE�o�oro�o�P(�Qϳ_�h�o����<*u�U�N��,��3lC�FXfr��r��t��.3��}��|k����q'�3�JJ�}�y
��.��(R�@�{�P�P����ϭ� ���Ώ�����M�8�`��{]�l��q  fU ��H�џ���������`��L�:�p�^��v�0������ƫ)ZƯد  ( 5�'� ���<�*�`�N�����  2 E���ާ�E�L����ˍq��B�0�#��PC%��0��@�_���
��.�@�R�'������ϟϱ����ϧ�?)��ç��%���r}�v��
 �� ?�Q�c�u߇ߙ߽߫� ��������)��y����n{V{H���$PARAM_M�ENU ?�u��  �DEFPUL�S�l	WAIT�TMOUT��R�CV�� SH�ELL_WRK.�$CUR_STY�L�`��OPT����PTB����C���R_DECSN ��u� �B�T�f����� �������������,>gb�SSREL_ID  �u����vUSE_P�ROG %q�%8c�wCCR������y��_HOST7 !q�!���
T���9 �;u�_TIME���b�GDE�BUG� q�wGINP_FLMS�`̠�TR��PG�A� �|�+CyH��TYPEn�z�b\�/�/�/ �/�/?�/?"?K?F? X?j?�?�?�?�?�?�? �?�?#OO0OBOkOfO xO�O�O�O�O�O�O�O�__C_�WORD� ?	q�
 	�AO��bMD9 ?��bIM��c�TE\�c?X	��RCOL�e�Y�_Z@&L�  �p��`���d�TRACECTL 1��u�{� ���{ �� X Y���|���:d	fDT �Q��u_`$`D� � C��l`0 t� l`7asa�rboo�o�o �o�o�o�o�o�o# 5GYk}��� ������1�C� U�g�y���������ӏ ���	��-�?�Q�c� u���������ϟ�� ��)�;�M�_�q��� ������˯ݯ��� %�7�I�[�m������ ��ǿٿ����!�3��E�W�i�{�hb` ���` �Ĉ �����������������������_v�_ �T���_��_���ĥ����w�`~�`R��`�ð�����U����	��
��:�`"�` �ĳ� ����������1�C� U�g�yߋߝ߯����߀����	��-�?�Q� ������������� �"�4�F�X�Z�l�~� ���������������� "4FXj|� ������ 0BTfx��� ��ha���/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� �����/>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰ� ��������
��.�@� R�d�v߈ߚ߬߾��� ������*�<�N�`� r��������������&�8�J�\���$PGTRAC�ELEN ��!���c���x�_UP �������������x�_CFG ������.������� ����� ���{ �����DEF�SPD ����-�� �x�H_C�ONFIG �d�����!�! dnMȇ� -�qP��c��x�IN~��TRL ������8�PES�]�����m\��x�LID�������  LLB 1Ǿ]	 ��B&} B4M���!��f`��� <<7 ,�?��� ������-// E/c/I/[/}/�/�/�/�/�*y???K?��D?�?t?�?�?�	G�RP 1�2�G�  ���
�.�A�PH���@B��A} D�	� Ap	@�r�$I4Imm �`�?�PN´�CiORKB�@�A�O{O�O��O�O�O�B��B�C5	_B_T^>_ <�oyQY_�_U_ �_�_�_�_�_q_�_4o �_DojoUo@z�c�oc�
o�ooo�o�o�o >)bM�q�������b:)�c�)
V7.1�0beta1� @�{@�?�A&�H�1=��C� CzB�O�D71� e�C�� b�ߛ� D�w�A@� �1B M@�1C6�1 �� �!�!#C�����B��0L ���%���0CRL���	����AK�33AFff@s�33BZ�Z��!A��ffA�33@�����^�#E�N�������O ��Fq���m������
�KNOW_M  ���SV �]
���oQ� c�u�Ɵ������ϯ��,MM�3�] ��M�	����C���:�����Ic�$@>� y�u�X��� MR�3��eT�J����C�c�U����OADB�ANFWD� S�T�11 1ϧ��?�4EOAT� with to�te�B@?�  ��L�33F����G�3F���fc�]�no8f�Ms� ���� �Iش��������� ��/�a�S�eߪ߉� ���߿�������L�c�<�2G��4/� � �<��X��03 n����<�4��������<�5�&�8�J��<�6g�y�����<�7 ��������<�8X1C<�MA'�-D�k��OVLD � c3��>�P�ARNUM  �J��\�39�SCH�	 �
IW5�iUPD�dE|���_CMP_���� K�6�'3��E�R_CHK����3�����RS8ư*��1_MO'�J(�_7/_�_RES_GF��c
���/d= �/�/�/�/???I? <?m?`?�?�?�?�?��#m��,�/�?�%�� �?OO�#�3OROWO �#f�rO�O�O�#��O �O�O�# �O__�#�_ /_N_S_�"V 1��J�/���[p�M"THR_IN�Rư��3�d�VM�ASS�_ Z�WM�N�_cMON_QUEUE �J�X3�/�� _�N��U!Nf:hQcENqDVat/piEXEo�pe�BE~``oQcO�PTIO]g}+T`P�ROGRAM %4j%S`�_8Rb?TASK_I��nOCFG �4ox�([pDATA��]�d{@ǀ'/�� 2 u<Ya�p�q�wY�v�q�y�u�u�w�s��~�q � ) ;+ ��-��g�>�) (G�H�4�F�l��R��)�I � ����� ��Iۀ����I���Y���0�0��y:��ZqINFO��	ը}(��+0�B�T� f�x���������ҟ� ����,�>�P�b�t�������wI �֨| ��9ZqPK_^qq�dy �ۦENB� H����2�%�G^q�2�� X,{		!=���q�����$U�!������T֧_EDIT� �d߿�WtW�ERFL�h�S9�RGADJ �κAйp=�?zH��Q� �Ta��/�?�A�z���p� <��)%DIAG���Ϻ�	_¸��2�j��	HK`l���RBp>���UU@x��*z,�/.� **:7�P'�9�Yߺ�P>����@�u�ߴب�Yz�8>��:�߬��߸��ߺQ�PA�����g�%�7� L�v�����t�������r����>���v����A P
�^�X�j������� ������P��L60 B�f����( �$�>� zt� /���� �l//h/R/L/^/�/ �/�/�/�/�/D?�/@? *?$?6?�?Z?�?�?�? �?O�?OO�?O�O 2O�OnOhOzO�O�O�O�O�O�O�	w�_�xo_�_�T�t$ �_��[�_�_�_o-oZ�P?REF �j����
 �IORI�TY�gն�$�MP�DSP�a����gU�TFv��ODUC-TCqκ0o��;OG��_TG�Hr�Һ�bHIBIT_�DO�{TOEN�T 1�λ (�!AF_INE��`epw!tc�Љ�{!ud���~!icmX�]��bXYc��μ;�ya)� D�$�6����_�B�N� ��r��������̏	� ��-�?�&�c�J�����I*�cc��j���%G_xݟ�yb>�%�"օD�/N�˟@�����������,  �``Ρ���������
e�0�Z0����#��5����ENHA?NCE 㺝��AЫd/���|��fId��Qocc�$�PO�RT_NUM�c��e$�_CA/RTRE{�	�ZSKSTA�g2{S�LGSbp�	����Ú`Unothing��zόϞ��7k>�TEMP ���i��#�b�_a_seibano � o�C�.�g�Rߋ� v߯ߚ��߾���	��� -��Q�<�u�`��� �����������;� &�8�q�\��������� ��������7"[ Fj�����|���VERSI�`��g. di�sable����S�AVE ��j	�2670H72%2��!������ 	��bA_+/�ce,/U/g/y/�/�*D,��/˭�K_p 1�	��w ��:�
W?+?WB`URG�ET�Bp+~�qWF W0'q�dj��fW^px4��a��WRUP_DELAY ���k5R_HOT �%fV�a���?�5R_?NORMAL�8�bx�?<OGSEMIO�AO�O@aQSKIP�#���3x��O� �O�O_�M^]<_lS@_ f_x_�_P_�_�_�_�_ �_�_�_,ooPoboto :o�o�o�o�o�o�o�o :L^$6� ����� ����6�H�Z�K3RA����Kh�H��t�_PA�RAM�A2�K; @g�@`�&j�W2Cu��BÁ�C�&ձBt�BT�IFy4�RCVT�MOU&����t�DCR�#�I� ��AE���_E7�iE�e�7D�C��ϚB���Hš���� ]�������� ó?2O��Ҋ�O���_ ;�x5;���0;�i;��du;�t�<!��ذ���&���J�\�n����������ȯگ������R�DIO_TYPE�  �-��EDV��T_x����X��BH�#E��j����nz� ��B�� ��Ϻ�������=� (�пn�mO��$_��� ���������4�"�X� Bׄω��P߲ߠ��� ������
���T�v� {�ߜ�6�������� ����>�`�e���6� ��2����������� :\�a��B� ���� �$F K]~��� ���� /BG/f (/z/h/�/�/�/�/�/��/�/,/R/C?�j�I�NT 2��9���4�G;� �?�;�x ��?-�f�0 �? �;?O�/OO/OeO SO�OoO�O�O�O�O�O _�O�O=_+_a_O_�_ �_}_�_�_�_�_oo �_9o'o]oKo�o�oyo �o�o�o�o�o�o5�#Yf�EFPOS�1 1�9� � xAT HGOME��Ճ��(�1���z��lu��
�Ż�����x�����(�=�5�}@N���=1?����?�H�3�l��ABO�VE LEFT JACKP(�Ň���+^��H�~�F�f#���4���+�ɏ���|�~���ڍ@���z���RIG�H����,^�@I����G�*;��"y��nʿ�ʏ܏� �"�\���X�џl��������+��O��E�O�pchangeO pos�w�g���?��x=�̅��<<!H����%?�N�p�����MAf0� 1��d��ɾ�I�/���E��<Lu'����������ί��2��e����>g�࿊H��<ǘ���x4���"�8�F���3c��f��ʣ���
ٿ5S��;j{�?3k����������At Palle?t Stop餡��o����>�����=�9)�D��t7>[����(�6�H�a���p����ҽվQ@����8xv�տ�T[��^���ϠϮ���ٴ��q���d��>	�
��
Ee�b����謹�����&�8� 4|�r�&��=������6K�f����"�4�^�zߐߞ߰� 㡉s����69�Յe�����4"���_b��!����'�p 6|�t���B�D=�E���	�I�	oK���/���Fc j�����<�M�8� q����0��������� ����7��[m T�P�t�� 3W�{� :��p��/� A/�e/ /o/�/�/�/ Z/�/~/?�/+?=?�/ �/$?�? ?�?D?�?h? �?O�?'O�?KO�?oO 
O�O�O@ORO�O�O�O _�O5_�O?_k_V_�_<*U}u2 1�3_ E__�_�_!o'_Eo�_ ioofo�o:o�o^o�o �o�o�o�oeP �$�H�l�� �+��O��s�� � 2�l�͏��񏌏��� 9�ԏ6�o�
���.��� R�۟v�����ԟ5� � Y���}����<���ׯ r��������C�ޯ� �<�������\�忀� 	Ϥ��?�ڿc����� "ϫ�F�X�jϤ���� )���M���q��nߧ� B���f��ߊ����� ���m�X��,��P� ��t������3���W� ��{��(�:�t����� ������A��>w �6�Z�~� ��=(a��  �D��z/�'/ �K/��
/D/�/�/ �/d/�/�/?�/?G? �/k??�?*?�?�_�T3 1��_`?r?�? *OONOT?rOO�O1O �O�OgO�O�O_�O8_ �O�O�O1_�_}_�_Q_ �_u_�_�_�_4o�_Xo �_|oo�o;oMo_o�o �o�o�oB�of c�7�[�� ����b�M���!� ��E�Ώi�ˏ���(� ÏL��p���/�i� ʟ������6�џ 3�l����+���O�د s�����ѯ2��V�� z����9���Կo��� ��Ϸ�@�ۿ���9� �υϾ�Y���}�ߡ� �<���`��τ�ߨ� C�U�gߡ����&��� J���n�	�k��?��� c����������	� j�U���)���M���q� ����0��T��x %7q���� �>�;t��3�W��?�44 1��?���W/B/ {/��/:/�/^/�/�/ �/?�/A?�/e? ?? $?^?�?�?�?~?O�? +O�?(OaO�?�O O�O DO�OhOzO�O�O'__ K_�Oo_
_�_._�_�_ d_�_�_o�_5o�_�_ �_.o�ozo�oNo�oro �o�o�o1�oU�oy �8J\��� ��?��c��`��� 4���X��|������ ď��_�J������B� ˟f�ȟ���%���I� �m���,�f�ǯ�� 믆����3�ί0�i� ���(���L�տp��� ��ο/��S��w�� ��6Ϙ���l��ϐ�� ��=�������6ߗ߂� ��V���z��� �9� ��]��߁���@�R� d������#���G��� k��h���<���`������A��*S�YSTEM*��V�9.10170 �G9/18/20�19 A � � 4��#51�_T   l �$COMMEN�T $EN�ABLED  �$ATPERC�H�DOUT_T�YPE� �IN�DX��	   w 	�TOL��HOME�  
i6qw���\�� Hi7q��*<N +�i8qq�p���� i�SMSKr � $MAXjE�N���4i MOTE_CFGr? T $�$"�" �#IO �*I�, �!LOCAL_�OP�%�#STAR�T{!��i POwWERr m /FLAG� �"�"�r , �&$�DSB_SIGN�AL�"�"UP_C�ND�!�S232��% � ���DEVICEU�S�#SPE �!P�ARITY*4OP�BITS�"FLO?WCONTRH �!�TIME �"CU��0M�"AUXTA�SK�"INTER�FACi4TATUf�0F A0CHr �	 t�OLD�_o0C_SW"F�REEFROMS�IZ "� GET_�DIR�	$UP?DT_MAP "� �Td ENB"EX�P0JC!`0FAU�L@EV!�RV�_DATA�1
 � $d@E�1 �  ? VALU�yA> `FGRP_ ��"dA  2
� �SC�"	�� �$ITP_�vB $NUM�@OU�!�CTOT�_AX�1�CDSP��FJOGLI�3F?INE_PCZ1�1OND�Eo!�@�6=K+@_MIR�ATmP� TN5XAPI >0!RE_EXXP2D`�A5 .Q�"�APGmV�BRKH�11FNC:�@I:!  �R#�R�BP!@D�!�C1POBSOC�F� N�U�DUMMY163��BSV_CODE��!*3FSPD_O�VR |@�LDLb	SORg N bfF�P2g�@OV�E;SFJjRUNMc!!�SFff�!SUFR�A|jTO�4LCH�DLYWRECO1Vd �@WS @�P��e�@RO�3�QP_~f`   @� �Su@NVE� !O�FS�`C�@ "FWD.a�d*a�Q�QU�P�TR)1o!_VQF�DOQVMB_CMt�!<pB�@BL_c (S^rdq2ncV�1 "�@s@�CFbG_wrXA�MpSRp�0�u�b�_�Mvp�2M�@�"�`T�$CA�@�pD�R��pHBK!A0F�I�O%��!"�PPA	�5��E�-��u�"��bDVC_DBG  #w�1A2w��b�!���1���s��3���`ATIO� �1�0aqU #�@�&CAB P " "P�d1 �x!!�@�_�00FSUBCPyU2PSIN_0Hs�t"@1D�ws�t�"~�Q$HW_Cq  �0S�$�|�wq
 @~|@�$UNIT�T�����ATTRIx3@��PCYCL#�NECAۂBSFLTR_2_FI-#�/9�"6!!LP[CwHK_�0SCT4SF_��F_��.����FS!1�r��CHA�=��o�r�2n�RS�D�`2�Q;C1� _T�xPROǀ6s�0KEM _�@�ST\��S�|@\�wp�DI�AG1ERAILAiC��*�M�@LO�P4!�V4�BPS�B"� #���sPRx�S&$@ �M�Cj�\0�	�cFUNC�R~�1RINS_T$A0 ��m��1RA~��@�; �p��p �t��W�ARBP�CBLCUR��ǴA����ø��DA�P���ǳ��LD@�P"�)��A��.�)�TI:�IſA�|@$CE_RIYA�1+2AF:�P91�t��`z�T2�C�/C��qqOI��9vD�F_Ly ~bA�0L�M�sFA�`HRD�YOBQ�`RG.�H���4Q 	���MUL�SE��3CI��P���$JjJ,bAg<kF�AN_ALMLV�)3H�WRNO�HA#RD !F�P�2��!2Gф1�A�U_�`0F�AU�0Ra��2TO_SBR�%���@���l�u���MPIN�F�`�������REG&NV@��V5D� NHtFL}��R$Mʰ��3I��p�|@V�]�CMj�NFƑ !��?ppr�k $-!$Y���A �B�As o� �eSEG���C�P��AR�@�#�U�2�S���rUAXE��GROB�JRED&�FWR�`�Q_#��SCSY�P��PE�SO��WRI�`��{�ST�0�C�0�P `E�� ? ��)����@B���ar��5��pOTO�9? �`ARY�C��0�˄="�0FI{P�3�$LINK��GkTH��8@T_����a��6�BXY�Z!B
7-OFF��`����B�@b�r�a)0@sFIʐ��0*3�Tb��D_JZ1|Bb��"��Х���8�Bg0������C�!bUDUt	r��9*�TURJ�!XP�4����X^��p�FL �`����R�6��30�Bq +1? K PM0D�U�3S�-�I�:�I�	CORQ���A���wq-�xPOA�z!b�$3C�A��$OVE!��M �0!��8%��8%��7&��16'$A6'@5$AN s���8!z���!/Pw  ��!0%!<'�%���%L\#�AERQ��	.�!E�`d@:��$A�!|@����������AX�c|B������� Y5�e9�e9)�d:�� d:, d:K d:� d:+d:1�d6��a9��q9 ���9���9���9���9 ���9���9���9�1�9oDEBUs�$n�`z�⢢ArAB���.a#V�pr� 
�B�����Ewq�G�Q �G)��G���G,�GK �G��G+�� z���.sLAB��o��|�GRO���s��pB_ȡ�&{�ã� ��КV�Q��U���VAND�.��$��!��g �q{��'h��6h� NTZмcY`VELΡ�$ca�kf?�SERVEY`�� $����A�!�`PO�bs�Ap���a�b�!�� � $�bTRQ"��
�c.��`�gz��2�fX��_ � lX��q�ERR��q�I�pg`�$,qTOQ�$� L�c4k�?v��G�e%���cRE
� � ,�a�e�`�"RA~�q 2 d�r�-�|t�` ���$, ͢��S2 ̩�aOC���p � {COUN�T���`��FZN_wCFG�a 4x���T�p���CsМ@�q������ ��@M=�!Ҡ�`Հ�#5!=�u�FAg��%u�y�X�u�UqH���d��P��Ω�HEL7��� 5� B_B;AS�RSR�V�E�S��B��1hw��2*�3*�4*�5**�6*�7*�8hw���ROO�op�� NL��AB�c ���ACK�FIN�pT�!�M�U����a���_cPUt��OU�cP~���ivb�}�?6�TPFWD_KA1R1q#� pRE�d��qP���s�QUE�@�� ltЇ�IKЀ�C� �h`�SCEM�A���A��Aq�7STYɔSO����DIՑ{�7�u�>7���_TM/�MANR�Q� END���$KEYSWIT�CH�-��~�HE�BEATM`�PE��LE0r�Q�P^��U,�F��-�S�D_O_HOMx�Op�6��EF� PRx9�(0�|�֕Cx�O��p�qOV_M�s�Y�IOCM���A�`��`�HK�� DH�G�Urs�M��xG�X FORC �7WAR�� �p��OM��  @��D���U��P��1(z�]�|�3z�4���*�pO=�L`��r�OUNLO�t�ěED��  �p�PHwDDN�a �`�BLOB  ^��SNPX_AS�� 0D�ADD|G�I�$SIZuq�$VA�PjuMU/LTIP�����A`� � A$�Ь�� ��S7��QC,py�FRIF����pS]�oɰ�i�N=F	�ODBU^�8`�zսӸ٥fw� �IA`N�������S�>�� � #�Ir�TEm��SGL1�T��^&)�J�S<G�2�STMTkc�P��o�BW 3�S�HOWk���BANw�TPU �+��h��P�V� _GY�;  � $PC�P�p��#U1FB\�P��S�P��AԐ��pVD���X�!� �qA00d1��9�@��9���9���9�57�U67�77�87�97�A7�B7�n�9�mQ:���9�F7��0��C��Р��]����w�1��1���1��1��1��1���1��1��1��1���26�2C�2P�2�]�2j�2w�2��2���2��2��2��2���2��2��2��2
��36�3C���]�U3j�3w�3��3��U3��3��3��3��U3��3��3��3��U46�4C�4P�4]�U4j�4w�4��4��U4��4��4��4��U4��4��4��4��U56�5C�5P�5]�U5j�5w�5��5��U5��5��5��5��U5��5��5��5��U66�6C�6P�6]�U6j�6w�6��6��U6��6��6��6��U6��6��6��6��U76�7C�7P�7=IU7JI7WI7dI7qIU7��7��7��7��U7��7��7��7���C�VP\�U�b"��¶P�
�Ҏa#� x $TOR f������r�`R�`ڀ�TQ_�pR�`Au�a�8�ndSmC��e�5f_U��@a�YS�Lfp�`$ �  #���$���ג�� ��<ld��VALU$�ߐ�2�a�hF]aID_YL���eHI�jIN�?$FILE_��df#�$��XfSA�q�% h�P$pE_BLCK`�1rL�:xD_CPUJy$�Jy �/��ot�pY1� ��R & � �PW�p�����qLA�q�S�p�t�q�tR?UN_FLG�u�t �q�t0��u�q�t�q�u�H ��t��t  w�T22�_LI`��'  ��G_�O��:�P_EDaI��0���:�(B��ɲ�Eqk�,��TB{C2#�) �(�`$��p����:�FT��\��ãTDC�pA���Q�ɀM�PÆفT�H�Ѐ���S��Rx�����ERVE����ã�ፂ� *X -$H�LEN��U�ãH��cRA\���\`W_a�ws1H��d2��MO$Bq��S��ҐI�1b`�a���TH�̛DEܕ���LACE�cCqC��1bp�_MA	�pۖ���TCV�=��T�>�]�S��ړ���JΠA�M����J��!�ڕ)ǡ�T�2������ٓ��JK�V�K\�� �����J����	�JJ�JJ�AAL	�?��?��9��=�5��p�N1�d�p�/��dL��_x_���^�BCCF��+ `�PGROUP�`M����N��Ca�~��REQUIR��ƠEBUx�D���$Tܐ2*�E��8��Д�, \B`t�oAPPR��CLb�
$K�N>�CLOD��N�S�c�ڕ
��.L�- ���M׀�8o���_MG�Ѩ��C#�%p�ȧ����B{RK��NOLD����RTMO9�������J9���PA����������]���f���6�.�7.�?���|C���.� ���o�\��� ��PATH�ױѧӱ�t������-3a��SCA�x���?§�ING�U�C�����C�UM�Y��vp����a�#�2��2�H�2�PA�YLOA��J2L��PR_ANρs�L��p}�y�m���R_?F2LSHR���LO~�U������ACRL_:q���� �e�g�H�`b$yH��%�FLEXA�u��J��/ P+�����.���@�G�0 :T�f�됷����i�h��r�����F1��0����ɟ۟���`E	��-�?� Q�c�u�����7T�� ���D f��̯ޯ���T�5X=a>� ����%���,� >�B�K�9�]�f�x���朹C_A�1 ������ο࿄`�PATI󱥠EL� ��3j��J�0�JE��gCTR �DTN�Q�6�HAND_V�BbA�`��2 M$�F2����c�SWA 	����3?� $$M���� �P���8���<� �5��6A�`j���aI��QA�̖`��A��A��P@��cp��D��D��eP��G�p�IST��h�A�ɼAN��DY�p <����4&E��I����� ����l�������P6�?�H�Q�Z�c�l��u� ���4 �0���� q�Up���QASYM��<������3"a������_ �����	�d�8)�;�M�_�q�Jx�)Њ�p�c�i��V_VIr3��hp��`V_UN Y��`s.#��J��%r SU%r��)t��6tZv�퀥���)�
���u��2�:��1���HR��w�5�2�qT�N�DI���O�tv2�pN��6 > -BIaA-���'�J 5c5�M ���� �p 7 �[ �1ME�� hP��r7aT�pPT�` � ��x����$S�o`�}�����T�`�� �$DUMMY1�H�$PS_G RMF	   ��ӆ��7FLA��YP�����$GLB_T �0�u�x�\��� H1�T�8 X+�뷂�SuT���SBR���M21_V��T$_SV_ER��Ob`LN�f�CL"�N�A� �O*��pGL�`EWβ�9 4����$Y"Z"W��頲ᒜ3AQ������U.��: �Nː�`�$GIX0}$�� 9|Г�ʐ���; L���ab}�$FabE��NEA�R� NNF;�� T�ANCNv1JOG���� <�0$JOINT�� w1ޓ�MSET��= E �E!�K� S�"����!��>� �E U�?��LOCK_FO��1�poBGLVK3GL�TEST_XMA�N��EMPw���	� �Р$U�� #2:�ʓ/�;���04ՠ/�9P�CE�����P� $KAR�M>�sTPDRA��m��d�VEC��~�h�I�U/�<4�HEנT�OOL��VR�E��IS3��ò6�Q�D ACH���=���O�Ѐ�3>!���SI1�  @�$RAIL_BO�XE�s�ROB�O �?�s�HOW�WAR-��Ѐ�ROLMۂEū!�V�p�!�8 ��O_F� �!s�HTML5��q �>�ݱ��?�p��R��O��@`�� y�}���OU��'A d��+�97a!2|�!Р$PIP�N����ݱV /���~��CORDEDՠ��п�8�XT��)��p� O7� B 7D �OBSA%3 ՠ^�MѼ��M�a`'1wSYSM�ADR&1��px�TCH�0 7C ,�EN�r]�Aܡ_��Դ!A{RD�pVWVAS�?D � s�����uPREV_RT~`Q$EDIT��_VSHWR�!:�(�����`Db����5�.!$HEA�Dra�pO��a�K�E����CPSPD�f�JMPj�L�uCg�TR� �EU�TR��I
�S&2Cl0�NE��'1b7TIC�K�aM[�v2��H=N0�F @WЭ��%n�_GP���^�gSTY���LO"��������G tk 
��G��%$����=:�S !$@q g��$��P�P��SQUg���a�TERC|�!G�S�$H �F��' ��'g��C O}�p�FR IZ����ρ�PR3�܁����P9Uq+_DO@����XS��K�vAXI4J i�4�UR� �@'2&���x֗1� _����ET�Pޢf��U%I�F�WJ�A�A�QÄ9�>0 ���{SR4Il�� �9"�:�6�2 GIILAGL QGLaF^x�I^�$�R|C��C�Zo�lo~o�d��SC
� oJ hs�DS��n�SP!�x%AT�O@�2,��⿂A_DDRES��B
��SHIF�#&�_2+CH&0t�I)��!��TU)�I�1 }K��CUSTO�*&�V��I�L��򨨌!�P
	�
��V8��;U�M \����A�I�<���W2C�C���):��l�W1�T�XSCREEO�Nz�pe�TINA��x���4�����sQ_�"�PO T�� i���h�E��6X��8X�4�RRO*PU�`��`��1p`�UE��GP ��P���S��N��RSM��NU<�0���vaA�pS_ē�F@cqA�I�Gc�Cʢ�]B�4 2O�0U�E�TQ�y��F G+MTmpLGqgU�yOz�&�BBL_�9W��U�R �I�!R5O��-RLE�"8Sx%��"7TRIGHAS�BRD{��!CKG�R��iUT=�hWeQWIDTH�+�o ��큭��@Ix�EY� T�S��D�-��=BACK+�ۂ4�U�[�FO*��W�LAB6?([�I<�΢$UR+�`��0�Pa�HA T 8�qU�_N��"?bb�R��Т��ˁ�AR-`O�!U�U�����bPUMP�cRޢP�L�UM�co� ERVH�����PP?��TVY�� GE b&�� C�&W�LP�e�E��=!)�g\�
x]!
xװ	yU5{6{7{8�b���p� ?�k4��ױ�ȡS��U�QUS=R��W <��a�1U��#�FO� �PRI�m��{q�p�TRIP	�m��UNDO�X� n��pP7�O�`'�� ��� Y:b�pG V�Ti�+!�!5�OS��J�R� B!���1�Z������q��$�A'�U�a1�[z���p�C�b�!�OFF���2�\6���O � G1Zs���[s�GU��P�{�-�(!7��QSUB򂐰�RTs��]��T�u����OR�}�RAUD� ~�T����c�_��Ε�^ |��OW�N$���$SRC�(@�@l�D����M�PFI$�S!� ESP'���0���c<�g�ɲ�p����A_ `&ÀWO2�����7COṔ$� &��_���w���~�WA
�C���[�1�Z�ɲp�p��C�1 `�2?SHADOWl ��~͡_UNSCA��8ͣ�TڣDGD�eяEGACq�7� P�PG�2a:bhSTE4Q:�Ox`�d�kPE�bgVW��62RG� �Ab y���0�MOVE(C��ANG�D��؃�������LIM_X ̃��҃����ı���C`K��p� ����VFi �~�B�VCCM��c�2C^�RAO�@�z�\� 5�NFA���Z�E�a�pG� fAPb��&�DE^��
1�.E��Ad�# ��z�Dű�Ȏ�dcpC���DRI����j�V������� D�tMY_UBY�tE�q�z�)A���0b<�@ر�O�P_㠴$�a�L1BM4Q�$��DEY��EXXP5C��MU��X7����v@US��v �p_AR�1���p� ��G�PACI�g�󑋴���؃�җ��ҩC��R!ETb�!q�:�����N��e � i�Gk��P�29���Ra���f �P�`A�Q]�	v�H�R6�SW���$�� O�q�QA� ��EzpU<�]������HKA�g�`��ꏱ� ���0��EA�N��Z�A`��a���MwRCV�Ah ��`UO5�MA`C�3	=�8�6�=�REFW_� F�1񵲸��pB���@S���d���F���_� �����4�4D2���0#�/�.�Di ��H�l0z�#�q�$GROUv ��0�mdE�w�dO�,!2e�@0�0m08�Pf�#,!X�R@� UL��g6��CаUah�Д NT1�����na��q�� LK�
[�
na��q1�T�DDj� tÀMDi�AP�_HUZ���VSA.��CMP(@F\um]_t!R�S!�d�X���GF�����k� �`M8�pAP0�UF_&@v�/��uROKP�2��7դ`F��P��URE��RA&��RI��_I � g��������ȹ�,҃�IN��HT$#��PV��ײ?��#{S�%W��'熡�Á���-9��LO�����#P9��\1uqNSI�VIsA_Z��0l �+P�HDR �P$�JOupR�$�Z_UP԰-BZ_LOW�5y1�GaRӰ[AL P�W�B��1y1- \@�g�0@�þ�m� 0�P�A�Q �CACHc4P1(EO1��DI�aT���CӱI�F�1�pET<PoF'$HOA`ܒ-@��öb" �FP�R����aT��VP3�.��B_SI	ZZ��DZg��H�1�G̖�|SMPZg�IM5G[�N0ADMYw��MRESmRWGP�M��ND����AS�YNBUF��VR�TD�U�TQ�COLE_2D״�U2܀%C�U��[@Q���U�ECCU&�VEM��(EbnGVIRC�MQ�U�S�b�Q&0LA`+���(��<�AG�YR��XYZ� ���сWj�h�!~dS�,`TE���IMea�VGb�cEGRABBn�YR7� E>n����CKLAS*@��A�K@o  �`T$4�p@��ܔ$As��p �v!��0b�#LuT�����7��r#��Ist'�Kf��BG_�LEVE����PK���Mf�PGI<pNaO7���i�8qHO�>��q � w�_�� �P�vS�0���R=O��ACCE��.�#�VR_c��M`$�؇����pARE�PA貀S�� Dq�REM�_B�d 0�x�J�MP  ��rt��$SS���d�0G|zQ@s  N2�SoPJ6NڄpLEX=vtȢ����� �DDR��$��Ӡh�}�\�4rP2F�u� i!?�V|_�MV_PI�S�u�T��z���j ��F�0�Z������y��!0���!��h�GAɕ���LOO~���JCB���~w�C���@֣PLCANҲqB�r�F"S O���P\�MQ�)�Ń���S+К�P��� �!P�nB�!��PâT9?��PRKE�N��VANC���R_9O�@v (B����ɳ�S��S��bR_}A�� w 4R��!�ΰ�p��k�x� h�ࢉ}1�W�OFF��v�F\`eD�EAj�
�P�PSK�sDM���� w ����@'�ry < ��-��UMMY�2�D2�M�'�CUS��U���z $� TIT>�$PR�+�3OPG�t3SFD�\�E{p���P&�SMO�|Ђ�K�YJ;����0Q_�E�}ЂX���0��@�XS�~ x>�0MSPD_���1ҫ`P�`�S40NB^�2LNTK3�M�>4�p�C�0#���1����'$��XVR&��bX�T6���oZABC=�K����-~�
m�7ZIP��Ђ�p�LV�CLw�~� ��ZMPCF��Ղ~���3�V�D�MY_LNϰı���� �ԃ �$�A ��CMCM�^ C�CCART_�G��P8� $Je�_�D�Ak�|� u� �� _�R�Y�z���UX�a
�UXEUL��ap���������������d�FTF��k�%�m������C ��w֟�?�Y�0�D�` � 8 �$R[PU2��EgIGH�X�?(� �����??�>� a��pf�q!6�$B� x�0}2SHIF����RV=�F����		$��6�C�0`�U�f�0�
Ks&�MD6TRb �V�Q�B>�SPHB�K�� ,� z��������0F� 5 1 �����  x�I t���	 � �� ��g R�&�J�n� 	/�-/�Q/�u/�/ "/4/n/�/�/�/�/? �/;?�/8?q??�?0? �?T?�?�?�?�?�?7O "O[O�?OO�O>O�O �OtO�O�O!_�OE_W_ �O_>_�_�_�_^_�_ �_o�_oAo�_eo o �o$o�o�oZolo�o �o+�oO�osp �D�h���'� ���o�Z���.��� R�ۏv�؏���5�Џ Y��}���*�<�v�ן �������C�ޟ@� y����8���\���� ����ޯ?�*�c����� "���F����|�Ϡ� )�ĿM�_����Fϧ� ����f��ϊ�߮�� I���m�ߑ�,ߵ��� b�t߮����3���W���{��x���6 1�S�e��� �A�G�e� ���$��� ��Z���~���+�� ����$�p�D� h���'�K� o
�.@R�� �/�5/�Y/�V/ �/*/�/N/�/r/�/�/ �/�/�/U?@?y??�? 8?�?\?�?�?�?O�? ?O�?cO�?O"O\O�O �O�O|O_�O)_�O&_ __�O�__�_B_�_f_ x_�_�_%ooIo�_mo o�o,o�o�obo�o�o �o3�o�o�o,� x�L�p��� /��S��w����6� H�Z����������=� ؏a���^���2���V� ߟz��������]� H������@�ɯd�Ư ����#���G��k�� �*�d�ſ��鿄�� ��1�̿.�g�ϋ�&���J��Ϲ���7 1��ϒ���J�5�n� tϒ�-߶�Q߳��߇� ��4���X����� Q�����q����� ���T���x����7� ��[�m����> ��b���!��W �{�(��� !�m�A�e� ��$/�H/�l// �/+/=/O/�/�/�/? �/2?�/V?�/S?�?'? �?K?�?o?�?�?�?�? �?RO=OvOO�O5O�O YO�O�O�O_�O<_�O `_�O__Y_�_�_�_ y_o�_&o�_#o\o�_ �oo�o?o�ocouo�o �o"F�oj� )��_���� 0����)���u��� I�ҏm������,�Ǐ P��t����3�E�W� ���ݟ���:�՟^� ��[���/���S�ܯw�x �����8 1� ������w�b������� Z��~��ϴ�=�ؿ a����� �2�D�~��� ��ߞ�'���K���H� ��ߥ�@���d��߈� �߬���G�2�k��� *��N�������� 1���U�����N��� ����n������� Q��u�4�X j|�;�_ ����T�x /�%/���// j/�/>/�/b/�/�/�/ !?�/E?�/i??�?(? :?L?�?�?�?O�?/O �?SO�?PO�O$O�OHO �OlO�O�O�O�O�OO_ :_s__�_2_�_V_�_ �_�_o�_9o�_]o�_ 
ooVo�o�o�ovo�o �o#�o Y�o} �<�`r��� 
�C��g����&��� ��\�叀�	���-���%�MASK 1�0�'�q��Q�XNO  `�~����MOTE  �� � ҕ_CFG �ݞ
��PL_�RANGّ?�4����OWER �0�R�9�SM_D�RYPRG %�0��%ڏ��X�TA�RT J���U?ME_PROg�y����!�_EXEC_�ENB  ��5�GSPD͠��;$�TDB2�D��RMS�D�IA_O�PTION*���7��INGVE[RS������H�I_AIRPUR(� ժ��
�F�MT_Y�TE�ۛ9��OBOT_ISOLC������K�/NAME���˿o��_ORD_NUM� ?��R���H722  &��@����.A������� 4������Q�PC_TIMoEOUT*� xQ�oS232��1���C� LTE�ACH PEND�AN������ُ׀Mai�ntenance_ Cons��j���"��ӄNo Usezݶ�|���������"�O�6�NPO��� ����3�C7H_LР	7�#��	��p�!UD�1:��r�RX�VA3IL�����5��_SR  ������~�R_INT7VAL���5�V�����V_DATA_GRP 2����� D;�P %���!������� >,bP�t� �����( L:\�p��� ���� //H/6/ l/Z/�/~/�/�/�/�/ �/?�/2? ?V?D?f? h?z?�?�?�?�?�?�? O
O,ORO@OvOdO�O �O�O�O�O�O�O__ <_*_`_N_�_r_�_�_��_�_���$SAF�_DO_PULS�ڐ��o�4�a�PCA)NҚ�4�aF��"�"5}�C�րր
4a���ĵѵ�
Xa�� ���o�o�o �o�o�oyo 2DXVhc�o�r���rXaXad�x�q�q8͑Tesy @�� ����y� ������_ �p.�T���.�k�}�����T D����ŏ׏� ����1�C�U�g�y� ��������ӟ�?�I��y��2�D�	����i�;�oJ��i�pl��
�t��Di��qha~J�� � �g� i�ha`ePaӯ���	� �-�?�Q�c�u����� ����Ͽ����)� ;�M�_�qσϕϧϹ� ��������%�7�I�@[�m�ߑߣߨ��+� ��������&�8�J� \��u������� ������*�/�l�F�0)�������{����� ����������/ ASew���� ���+=O as������ �//'/9/K/��o/ �/�/�/�/�/�/�/�/ ?|�5?G?Y?k?}?�?`�?�?�?0�����p+��0�0�0�0�d`qOO+O=OOO ]GnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o`�o�o�o�o�g��� d'���o,>Pb t������� ��(�:�H�Q�\~�����q�w��M�	12345�678��h!B�!��e���pc � ��$�6� H�Z�l�~������� ˟ݟ���%�7�I� [�m��������ǯح ������1�C�U�g� y���������ӿ���8	��گBH,�T� f�xϊϜϮ������� ����,�>�P�b�t�߫;�j�ߪ߼� ��������(�:�L� ^�p��������D������ �2�D� V�h�z����������� ����
߯@Rd v������� *<N`r1 ������// &/8/J/\/n/�/�/�/ �/�/��/�/?"?4? F?X?j?|?�?�?�?�?@�?�?�?OO&D߆AOSO�/xO�O�O���CB�A��j  W ��h2�b��} �H
�G�/  	ĩB29O _�2_D_V_f\�ogL���1�@3 4 5 6f_�_�_�_�_o o&o8oJo\ono�o�o��o�o�o�o�o�o�^P!r('r-?Qcu �������� �)�;�M�_�q�����B�A g@h@Q�B<��� ��Q  �ɋ㏖�ƂQ>Qt  �@�����`�$SCR�_GRP 1�"X�"al� �� ��� ��E	 j��r���|� hA�������������άM��@�D�` D�@|]��'��ᛊ\R-20�00iC/125�L 567890�PX�PRC2�L g���
V0�5.00 ���� ��vS�H�B��r���@a���a��S�������ǩ	�J�*�<�N��`�h���H��r���v�ѥh�D��|��JOC3�:���>����;	B��8������\��X'����ܾ�����@q��hh��  @&/nD����?�XC2#�r�_���%��ܟIϟ�;ϴEհ��T�8ﲕBǙ��B�  B�33BƘ��ŗ¨Î��A�@�����Ď�@9���� ?��ǎ��@
��ˎ�F@ F�`5�=�4�a�L� ��pߕ߻ߦ������ ������.��+�=�O�B�]��ߣ���� ��������!��E�0� i�T���{_���͟�������
����@+�&�,����R���h12#34f�x�F7O��A���������Y�$� �Q�� �'5JVh7  �����
/�"A�ECLVL ; !��Ѣ��"!L_DEFAU�LT*$}����uP>#HOT�STRJ-�"!MIPOWERF) ��EV%%WFDO�K& V%!"RVENT 11!1!w#� L!DUM�_EIP/�(�j�!AF_INExJ ?4!FT�/>>?b?!a�z?�;��Q?�?!RP?C_MAIN�?�8q��?�?�3VIS�?��9��?FO!TP&9@PU=O�)d5O�O�!
PMON_POROXY�O�&e�O��OYB�O�-f�O*_!�RDM_SRV�+_�)g_v_!RȊ�_�(he_�_!
��0M�O�,i�_o!?RLSYNw�*o�5g8�_Zo!R3OS�/�l�4Io�o�!
CE[@MTC�OM�o�&k�o�o!=	�bCONS�o�'�l�o>!�bWA'SRCE_�&m-�;!�bUSB��(ny�u?�9S�� #�H��l�3���W����'RVICE_K�L ?%�+ (�%SVCPRG1����2���3+�0��4S�X��5{����6�����7˟П򀃤��9� �_H���� p������E���� m��򁕟�򁽟8� ��`������5� ���^�ؿ��� �� ��(��֯P����x� �&����N����v� �������ƿ@�B� ���҂�ُ뀋��� ���������@�+� d�O�������� �����*��<�`�K� ��o����������� ��&J5nY� }������ 4XjU�y� �����/0//�T/Ɗ_DEV ~�*�MC:\+�8n$GRP 2��%k �bx 	�� 
 ,� �  k �k $bk 0Ak �  \$��"�" f�$�!Bk �$�%\#�#I�$�&�'\'�#�a1�!%�$*89#�$a1 �5)19?1'3�9e;C7 �%}515�?�'j!)1�?�C7�(�%a1O  ]qO�4�!	:O�"�$�/_0�� �� �Jk )k 2>�#uk U�k lk +k 'k U&k D�(�$�k U�k *k k �$�%5A9YAf��)	?�#�&DeAY1�5AO   bD�A�!p_C7"41)9y_  .H�_?; �Y�!)5�_gO oC3�$�YW0�_0�k LBk -�D%ec�#�k ��k N�$Y1a5==,
k k "8e�M�! �A�QY19�?cC1e �og�5O�_eA�9\ �#�_�mymU)�y���$Z� �k rk �@:Y1��m_ b�I���m��������� Ǐ�������j�0Q�����"�_0~���k �@X25��"��� k @���C7Ak .^T�AoC7�!��!a1�_C7�T�UqG W������-�����������{�T��z"k G�?0�k K&Dť�oC7f�Q���a�Q M�ݿKi���15�Q )�?;)1�Q)1i���# �9�_C7�%a1E_�Q!ҿ`���?��c�J� �ߙ߀߽ߤ������� ���;�"�4�q�X�� |����"�������%� �I�0�Y��f����� ����������!3 W>{b��h� ���/(e L�p������// /=/I(d ��T�I6 2�d@�@ԋ����@�t���n��%3=��G�I*g @#x���M�e@�F=�A��V@����?���-B^�:A���� �@�D{ϲB�k��*�^�8��x�'B����]���������I)%�GRIPPER�_OPEN _P�ALLET_RI�GHTI,T�O�a ��"H�B��`Aq�=�WJAs+�B�j���V5��"�s@�@�Ai�,?����@�p���O��V=A�4��c�;@�y��j��Q¾��C���V=?�B`�5�&ȿO�l��%*�R2s�4�� V9%PLA�CE_�0STIC|?I'T�Qbb%�?����f��@���@6���|k��/�V=�!���@�����T�h>�pA�������>V=B�*����s���������JB�ꗦ>� ��.��BE�Bd*+���_�AJ�X�?�?�? �@�b&�̖����@�IJ�=� ��g<�D�M*N�lk'� �@��bo@�i���>���RN��	K���`�����9j���mB\V>�tq��?�B��ͦ��?A�>�A�ǢJ�; �O(9Tb%>�m���������������}�M��V>���ʔ���畱A��A]	ƿ�*N�������X�>A	��Uu[��7Q*N��S�B��Ez�1�,�p@�k��J�CLAMP_C�LOSE���TLE�F�] T�	��b%�hΨ����>��=�:�������V==������ք@�J�A��A�A�%>��0�_ު����o�H>@����Uɰ��6��^@�Z�"�Bo�s��+�i�ԳA	7��Jo\fMING �_|eS�VH-����,��4[���7��VU･�4V>��@5�?�,^�@��QA����A%�tV=����B��.��ڶ�Ң�9Y�(C4V��~����·�"B������f��g����v_7mb�ko-3�3�b%;)�Pz�/�?��j�=��G���&˽��*Nu�5�O@?�X��@/Ơ��t]�:R�&_����#���r�����{��B�s�N_`P�[�B�$�����A��bAd����?B(��b%<���r�(��?��ъ=�D����}��$*NJ�$l����@�"�@K�h����b��t�B�����d�����Å�{��$B�+�>�U�U¨��B�r����z�A�Y)A�:�Ə؏��(���b%=�X��� iX?px��K�0�j��=����_����h�.?Q��߿�Z}�OO����|��^���8�@�[¿{��¾�)N���^���B������7A{��`h���ج��'���f֕����=����=2����߳��m;V=>������?��rSA�A8? ���o�f�G�o\8����,�gB������3����A��;�\e����}c�� 65>��G���.�O�@��g@��Ⱦ���9*N��
��(��B������(�ڼ@��RN�&A�V����������uL�B� a*F�OhL?�@+��&2	?���������Ep�O�O�� ��TČ�65�p�������B ���� �d�	ϖ��S�
R�e�?�)�����?AG�����x?�I�����2�r���B�q;yO�\?M�ڞ�<�b���> �@�KV��$ώ�KI+�,T�U�b%��N��1`@���꾎 �����=De�V=���Β��m�A�9�G�q�*Hk�«���%�=Ke�����@F����Z*Ne��/��sNB����A��!B,�x�A\q�z�T�_HE:�_CHE}C�T�W֖�ft���81��Q�꼌���ȅν`tVV>�A��d�7����Ap��ϑ�}��o	`�T������3��>@�1�U�G�`��T��RB�����G��A�qNA ��vB�\e6���ygŪ�b%@'=����:Amw=���:��[�?�.}>v2�:���� �6Z@԰W����z*���;����H��9���gJ	��BpN*N�{B�����B����By�zAN��B,h����f��@�Ƹ65�����>\d@0p��nq��K̻���V><���y�A��5@j��+@������V=C%&S?��f���?���ª��~��F���A�,b�;��C�.t@D/Ak�E�t�JAC�KPO7�8��@_T�ƹ�65=��9�B-�?��p����(A�p�@��*N����/�A���@z{�a�<��n-!�����B%b ������,��n�?��)8�*N�)��A�����!:��?G ?�3㏾��f�x��� ��TǨw&֬��u��X��^�� @����f��>�]R�*N�����L�'�������A;3ߊ@&��n�C��Aw���
�!�q���mߐA���~>�G����B���zA�<c��R|@��� ���@�K�b%�C.���t4�����@�jX��������V>���pǼ��|=?���A��J��ݔA�]%�[��p��؎��ΜB8�F��,@�~��B����?�g@�?<@����(�~^ �TȻ�65��!�	��W��B۾�CP ���@: y�n�;@��D3�%�:���^�AP���6Βʮ������)�r�H�>!�����PF�1��P��W�Y��@���h�7��c��*�PICK_INC�O9r*i�(T���������E��g�����Z�̨�"[m=���{�~dy@k��)@�@�5A P��}i�B@'B8v����@�u>��]�|B���RN1�������q����A��U����/����`��6�%���X��a-���̿R�<���"n��A�[��@�V!A��&@Q,^���ƾ2t�Bs�����#�@}����6bB�c�E�@P���m��B=ұ�� ������A!���/�/�O �T���~���#�@�Ҏ�At��E���;���m5�7�����y�AK;@�Kj�A@�����~�ГA��/��ݺ'�ry"��C2���~DK��A�(~��Y_����/@>2���v���?L����~�B��7�B!�[B�r�����>�+F�@B/Qn����56�A2���g��+���m�L%>-�Ћ����x�7�{�����¹eK��3��>.ٳ�A�9D���O?�R��?�1�>���{�2PAT�H�6/i�%T� ��&������@�(���~��D��R��ʮ��������AICm�*����"_{�Vr}Snߓ��Յ���@���,g½R�n���hL��'B|��/����AU���߰�F� ���63�B���?��)�M3���,DG�M��޺LV�@���P�K_����f�>�"^�{���J���Q@������T�2�"������B�	A�TM�B��A��o(o��� ���������??N��@�߿���OA�70@}��|;O���"�.�,���&���������@�����V������ÚB�_2�AR�A�؇A,����� /����;�p�����>z�&���-`����?7��>���4B�c�9���7A�zE='�*�����B����	�:�\���x�B�%Bi ����UB`@�����o�-=y���"�@���Z%�JOGG�1X� �?i����~�����>lL�������
?6��>�(�B�\�G���eQA��Js>�$0�� B�����:�����B��ZB ��A���:�@�+���e��%*��/@ ��*�آ1H_R�;բ�+��|>Y �?���K@~�
��ߕ�E��6~�ֿ���s�A;����_@D�v@���ڟq_�;�@���J(B���rB �}��_>.�
�A���i��@)���@� ��2A���6�uB�X��f������>O|��?�}�@~�T<U�w�θ�������A��D��@�U[@���׍��;�����*<B����B �b�3��&�t\A�B��z%�@%��|?#���0�ҿ<�yCJ�\�٢���_>Lk?��Y�@~�`���˧�E����$l��\A������@��>L@��VϞ�'�;�U���dB��eB ��s�>.&���A�����@w�e� ��O������W�ۢ��j>7�څ?�@~����\�E�k��?��:����VA�΀���@��D@��R�*߬0�< �����B���$B ����/>."*yAY�W�H�@j7����"��e�k�I�[�ݢ�E�g>.?�{�_@~���R��DU���W ��ʔ�A���%@��(�_�葹!�<7������B�o�BJ&R��d����A���@��ٿx;�Т�\��\���7�b>�!?�`�!@~B������E0-�?'0����A�[��h�@�#�@��8?���	�<�h����B��M!B���O>.#�B���!�@d\��B���,/�m�[��:���^>	��?���@}�޾1G��E �������Q�A���D�Ҹ @�U����<�������B��*qB7���D>.�SA�
�"��nѿX3��0A����F�,�2	=�$�<?�
�@}s�N�D���E ������Ċ�A����n��@��*@��z�u�<�����HB�8BU�e�^�@�A	hT��;�B��5���V��,����t��+��@|T��k�X�D B�����,��bo�����@�q�@�?�N��<�����kB���Bx���~�A*X���UU@��0��(\���(�<����=���{q�����D�=����T��A���O���Z}@��+�"/��=�^��QjB���nB����~�G�fѿ���fPj"���:�Y����(mV�����?�u@{��.���X�C:y��/� ��xA'�?���@�|�K����=����8�B��B?��%�7��
o��%1@��uX��:���:hcF?�j?�"	�ƾz�=�=�?�$�@z������!�CO��������% �A��A��S�R�@�,�?�;��=6�����B���B���9�v�~)Ζ����?w�U?�;O�%���=��@ �B@y}=�v���Cz�J����0��>^A������@�Ì��O���:��=J�����B�e�B%���~�+=�A`տ�D��@l+i��&p?�s)�O<�	_�+�f�?q~?��3�?�8)?n��+@����_�����Ƽ��A������&��@,BI^�����?o����B�i1�B `�Ed�~�*@�K����3@1�y�((\?����O�/�$�f�9��m�	���?`�1?���ֽ�����?H~�&��ss�A����9�@�2�@��������=����j�B��qB ��Y�ծ>x��q@Mڞ�R��@�o-?H?0>���o�o�z��"f���a
��?`��?ɛ���B���n���j8�A��}�?�@��@`�>��*�<������B�VvB ���<��1��P@E��|���^q> &p��%h�ߜߦ$�{Y��?_�c?�7�ｷ����4�!.�rq�%����6�Bi�q_����;����'��B���B ��{IJ���%�%@O������@��ڿ�%z�x��:v�_�(�f��a����
?b�N?��tc��ߎ������n�p�j�+�A����	��@�3�@[�I��k�:�{����B�R�B��\~�-E�@Kˡ>�>_p��!��;��_�3�E��zg?�g��?��Խ?�^ÿ�t�N*��necA��d��	ì��Q,^������9�j����B���B��~��m��@$����O�l@�PV�2˰>�)DCL���o�@��e*��H�?WE�?��E���y��i�B�T�q�����1@���@^�[Cj����8w�X��M�B�N��B/�s�!���{"Ғ�x=�ڒ�8�?O)E�M���@�#����|?^�}?ʰ�ؽ�Xk��T�#~�<�m��Aw�9��;|f��x����7a�����$B���B�B��.@�I|@G����������1s�?��ɥKPOۤ�_�E�%�e���������C���ʺ��[�'�=�񥒮N�c��fD3A��h��:R�@Ơs��VrSr^� y��6�i��l��B� >B�[�}�@3��?E���B��?�~��1C?���"���F�'����m<\�?����@z9���Q�A�'��Hbo��}ɲ���@���@��7 r^����7)6���B���FB���~��~@�*y@�&����#@�s�� ����߰6ߦ�[�A�*��VpM�?�@�?�#�?���@3��x���O�h�.2bcP�� ���@Oja�r^����9T����5B����B Y�<`�����Tp�W��<�b@/���;����
��$�
��",�Vurq�?��c?{V��?�k�@opﾄ�r^o� ���	 A��&����oZ�������:����(1B�8�A�+!�	��^�K��=C��?�=@b���3��M�+�E�.�Vxb��?�\�?oz9�?���@~kϾ��r^������7A����Ė��@`�@r^��C�<�����B���A����~��۶�'��R����v?��d�"&���ܲ�������"4�Ʀ�����+�������ҿX#X�=�Lޒ�E�u��qx�A��Z����������r^��!�;H����;�B�2��A��n���� ����_D>�_̿7���Ɔ���"8�e��#$6@7��@��[������`Z>��o���!���ΉcA��̾R�Z�1����~
�"��A�6����B��\BA��%��l��K��վ��>%*��@@Ca>�&OT���<��:]@6��@�`y���D���>�	��������A��ì�=ք@�ʔ��y�e����H)�F�.���xJB��]A����ǽ���@�T��O?+�{ޑ�@�O��O/E�A�z�9?UU�?��E/�%����DB~����l�ۦA�������@�K_@c��9�/o�Dc����E�B����A��g�~�&ꎤc**�k���@=Sv�"C=��=/ۯE�J���z?Y�?��[4�
�������B~D�v��m�A��������@���@�h0�?6�C�GU���B��J=A�'<�|��t����@7�5����V��*(�>�i{E��O*V̖��&�{?���@�����a�D@���������վA���F�c@��N��ZO3���C����u.B����A�۝��y����A.�v���@n7�' �� ??� �F�Q�e>����>�/������]�?Q�Z=��,�.^PK_���N�A����w����R������l�D������B���A�i��z�����` �Ș?�Z�m��#�?��)m~_?�?�bS�N�{п3�?k�qp?�mܾ��x��A[��=�qRE�A�zպV�@�P@v������HF�B�������B�lA?����y�K����ڞ�O�@9l!�P1�@&�Ro�Fե�_G�YN�� 8<?S��?��P1����� ��n�D@W@A��7���@��Cm@K��oH���A`������B��A�&���w�5��	���?��^��%��@j7���0�Yy�&��?>��\ʵ9+�' -?�SQ_?Ϭ��?N����z�v�d�A�`��� ��@� �@���a��@7����V�B��pZ��v��ꎒ���?s ��'E@���#�������_JH�n�ʺ%�?T]��?�e� ��Ͽ�!K�n�P�c�0�A�lk��Ew@߬�@t�T~�I@�?	�����~B����A��g�uR�����|�?�����]�3@��?��:,���5�Ut"�(F�?�L��?˞/� m
��K�V��D@g]qA�as�ٿ��@x�R�I�l�=���!�`B��A��߳�t2���{�?�p{�um��@l+i�$󄿋��4INT3�H&ş�V/1�>7=_�.���e2>��v�=��.������A?A�1n��W@�*�����oTF�>�����ZCB����A����t|�X��o A�I��D�?bi�1C� ̏ޏto´��V�2">6�8��'��j�\>?�4=M����!�% A�Y�Ͽ6Β� �����>�����O�B��A�ɥ��t�R��I|A��E�f��?z# �S@\�J��\��ؒ�>9����)>�֎?"���7���E���Q��}����<@�i�@�4+y��Ծ;��=����uMB��sdA�3��s7H2N��P���D����X?ֳ?o���	�����U�Zʒ�>���?!ﲽ^�9i�D	V]����>�dI�A��H�ܙG@�m�@�ˢ���[+����i�B���A�O.��r^�P��
=q#��B&!?���O�U�Z����k>�8�?���P}ƿ���V]<``�f���JB���@ο��@"��v�����;�*����9B�t*A�����p��V^����0=w @Կ�(\=��O��4M����6����V�>�Q-?�#�a�[�4���*o  �b��zA� ���?	�@�V��J���b�:~����AzB���A�����o�z��,@��s?��Y�@3�#�x�;�?��-ϻ�U���Ꙟ�>���?#g|�o�����0�_�^[CA���m��G�@ǿ��@�������9f������B�t�A���}�nx����.���?~�@1?�y�H0j�|��� ��Zʚ<>��?�?%�-�w1z�X���c��@�?��@Q�������8J5���$�B��XA�!���mI�F�X��B�I��u��)�R?���B�1CGKPOk�c�U��i���M�>���?#_�j�r�^2�g���A�t]�����@����ܱ���7*B��N�B�u�A�Y��l��q�x�@q��?DÅ贗������V1���>P������aJ>�*�<�c�.^,B����W�Aќ���AZ}���L�=_�.^��F�7��]��ugB����A�Bh�l�B�>��A�4��^k<=y�Ɓ�	���/�ؒ��V+�>9����'.��_��{>�`�<��$�.^-#���(Aק��C@��3J������n/��82	���[B�dIA�WM�lLr�����qA����g�?�o-�!���s)�/�?n��ؒ��V7l�>@��3�ҟ�b�7d>�R<���.^ǰ�����A�}۾?0�:�R����.^��7��8�L����BB���A�?hi�lU��N3�~���g��<�� ;��L8�?���;�/<��V8���>A^Z�#��t�a"~>�8��<�lF/X!s��A�x���ٿR�Z�mL�%.^�k��9����WTB�5�=A�~�l_�w�n�,@AT���`�]�� ��*H@?�9�������V;�H>H���%�g�=��1=0[h�^@����Ag �������P��Mi��^Л�9m`����2B���A����lh!���3�wP����=�_��2*�@��:_�?�O�ؒ���<ù����_�%>�?�Y=':?,4���.Br������^�����9�����B���A�����lr��_4����{S�>`f�@C���zo`���vV�:�G>Dp���}�he�>���=9���^�1����yA������Hb�o��P�^��Q��:<���<SB��q\A�����l~Z��PDx`���Z�m��:�@�UU�o�oؒ��
���d�>��I?(YO�O�>+��ʆ����h�kQ�A��J����X@ÿ��@ վ�o'�:�8�.@�B���A���k%�UB`���l���?��ž�1�?����R�?��R?
�? ��? J��?C �?�ӟ��Ihd�^�@�����A������,^�/Ơ@�U��z2�����:����|NB��p�A�gpj������P��0U@�0�1C��t�����֔�Ɔ���?"��?��?I/*?����Rmү�䠿��A�",��洳�W @Z��J�^��<�Hz��n)���A�y�j�`���x|0B����J�@?G ��<���05���|����=���4+��?D�W?����1�}����^��v�h���A�<���
�@��	@ec�j���:h����4XB�obA����i��@�@'P�%1�@?���&p>�%�2� oV�h��vV�J�>�_���k�_����?^�O=�x��d�7��p��A�>3࿺R��G��q�^�:H�;�N��R6B��31A�j��i��E.r�@�p{��B�?�п�3��>��n�(�f��R�f���?�d@�����
?�MJ��^>�ք���A���F���@��J@�������\�;H����B�v]A���e��r�����A�!�V���@fPj:���:�ڿT�h����z��?{�F�?s�R?�5��@����&���^�Ew�ţU�A�A�����@[�I�^Ď���=-���G�8B�D�A����f=x��İ������3?�?i� �.������d�$R�;:��?I��?�����K\��ڡ�^��c�xA���
��Ė@�7��
��Ś
�:�����B����A�A*�d{�Xr�G�?ǰ��R�&��%z��q�ߔߦ�h�%~	��4� ?@��?��⭾R�����oin>����f�"��P�@�zE@T�W�����9�������B�#�A񿃊�cb^��	���@�`��'E�@w�e�
!'�x�/V��2oh��'��:'�??���?�Ou�S��ȿ�����m���A�˞� ��?@�(�@tT���=�8[�����lB����A����b�����@5&�����7@d\����5�?�)m�*��z�h�2vV�~��>��i�z �ȿ��Y?dc�t<��1�s���A���>A���@��,2�R��9E����B��T�A�Z���bz�Z�^%%@>w��ke�[@N��GZN��<���h��5vV��>����q���Ƙ��?d�g=�x���B��>��������>\����d%�9�������B��A�Yp�b�Z��I|@� ��c��>ڬp�$��ֿ�d�7�y��;��?@[F?w޳x~��Z����P��`����H�@ǁq@i���þ��7������yB����A�	��`�����v��@	����p@Gȿ� �R��d�:�f�B�:?=_�?��r�T<�׿������e��uA����{�@���@lk�'*/���6�1�����B�S��A�Ns�_w����ϴ�@(���~@P���. ����d��@��KX?t���?oz9?ս�+@�Y��eg%2�����A��������԰W@n-$��^����8�����aB�ަ�A���_=S����@�%���?&�@3�#�((\~߈%�$W_�Y�F6 ����@���@��O�#	��K��B@t"Z���z��]qA��I�9�����*��Z������m"���L��B�R�B�`�¯I��$c*����]t�@�(?���"O�`?r?lR�$SE�RV_MAIL + v%HP��q2T�OUTPU� ?V��p@2TRoV 2f�  KP� (�s�  ���P"  �<_OVSAVE^\LY�TOP10 2�~Y d f� ��^B  �^@2�  �^@s�pT^@mQf��p�^@��pf�P�Q^@�r2c�P` &�Q Z�Vohozo�o�o�o�o �o�o�o
.@R dv������ ���*�<�N�`�r� ��������̏ޏ�����UYP�_NSFZN_CFG Z�KSu4mQ�U8��GRP 2����Q ,B   �A��v!D;� B}���  B4+S�RB21�VH7ELL;�Z��V���u:Y��u;%RSR�����F� 1�j�U���y������� �ӯ���0��T�u=�t�l��  ��Q%e�����s�s�w��"`�����@u7��	`�Pm����_HK 1��(b ÿ`�j�bόϵϰ��� ������
��E�@�R��dߍ߈ߚ߬ߨ�OM�M ���߬�FTOV_ENB=T��Q�U;�OW_RE�G_UI�ORIM?IOFWDL���Fx�V��P�WAIT�A�Z�x�XP<��T�u�TIM<���Ư�VA<P��P�_U�NIT����YLC�5�TRY<��U���MB_HDDNw 2~[ (` ��u5W�x��s��� ������������$�8�ON_ALIA�S ?e���Phe�QZl~��u6 V����); M_q���� ��//%/7/I/� m//�/�/N/�/�/�/ �/?�/3?E?W?i?{? &?�?�?�?�?�?�?O O/OAOSO�?wO�O�O �OXO�O�O�O__�O =_O_a_s_�_0_�_�_ �_�_�_�_o'o9oKo �_\o�o�o�o�obo�o �o�o#�oGYk }�:����� ��1�C�U� �y��� ������l����	�� -�؏Q�c�u�����D� ��ϟ�󟞟�)�;� M�_�
���������˯ v����%�7��[� m������N�ǿٿ� ����!�3�E�W�i�� �ϟϱ����π���� �/�A���e�w߉ߛ� F߬���������+� =�O�a�s����� �������'�9�K� ��o�������P����� ������5GYk�}'�$SMON�_DEFPROG &����� &*SYSTEM*���@+ �RECALL ?}�	� ( �}3x�copy fr:�\*.* vir�t:\tmpba�ck=>10.�$202.21:?19680 2;XM_o}4a�/8��� }�8s:orde�rfil.dat����J/\/n/}/mdb:�'/4 3/�/�/�/{�& �/I?[?m?�?#?� �?�?�?�/�/�/EO WOiO|/�/)O�/�O�O �O�/�?�?0?A_S_e_ x?�?_�?�_�_�_�? O�O,O=oOoaotO�O !o�O�o�o�o�O_�_ (_�oK]�o�_% 8��� oo�o�o G�Y�k�~o��o4�ŏ ׏��o��2C�U� g�z�����ӟ� �
���.�?�Q�c�v� ��#�����ϯ��� ��*�;�M�_�r����ਟ:�˿ݿp�xy�zrate 124 ������D�V�h��{��#�8:172�"�4��������� �ϡϳ�D�V�h�{��!��69.254�.14&�4:16120 %�7���������tpdisc 0�ߠҢߴ�E�W��i�|�tpconn 0�� �2�������z�:����=�O�a�t�1����� 6�������~�5��@�����K]��6��& :��p� �����I[m�� �6������� 4E/W/i/|//� �/�/�/��0A? S?e?x�%?��?�? �?�/�/,/=OOOaO t/�/O�/<O�O�O�L��$SNPX_A�SG 2����Q� � �B%��O6_ � ?��FPARAoM UQ� �	$[P�$r� 9X�T�P�POFT_KB_?CFG  �#U��COPIN_SI�M  [�R��_�_ocPRVN�ORDY_DO � �U�U#bQS�TP_DSB�^��Rgo�KSR �Y � & �PNS0001 �IONCHECK� T T_RIG�HTsi�$�ST�OP_ON_ER�R0o�B�aPTN �Up��A�bRING_P�RM�oBbVCNT?_GP 2 U�QPx 	�V�YeXP{�}n|��p�tfp��s�JVD7p�RP 1!^Y�P vqah����0� W�T�f�x��������� ҏ�����,�>�P� b�t������������ ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�o�l�~��� ����ƿؿ����5� 2�D�V�h�zόϞϰ� ��������
��.�@� R�d�v߈ߚ��߾��� ������*�<�N�`� ������������ ��&�M�J�\�n��� ������������ "4FXj|�� �����0 BTfx���� ���//,/>/e/�b/t/�/�/�/�/�rPRG_COUN�`�T�r�)ENB��%M3�T?_U�PD 1"�kT  
�/|Bd?v?�? �?�?�?�?�?�?OO AO<ONO`O�O�O�O�O �O�O�O�O__&_8_ a_\_n_�_�_�_�_�_ �_�_�_o9o4oFoXo �o|o�o�o�o�o�o�o 0YTfx �������� 1�,�>�P�y�t����� ����Ώ��	���(� Q�L�^�p��������� �ܟ� �)�$�6�H� q�l�~�������Ưد������,_INF�O 1#R5980Z�	 1�u��`�����  ������������\�������������h¤@t���~���� �D�^�@�C2�Խ������-B�&��8�� YSDEBU)G� S0�(�d;9c�SP_PASS�%�B?u�LOG �$O�\1  z(���?��(��.�  �71(�
MC:\�Ģ��)��o_MPC�� ��x��.���UD1���25��SAV �%��1���*��Q�SVb�TEM_TIME 1&���]0 0 a݆'�|m35 ������g'��z��MEMBK'  R571����x7�I�Y�X|80g� @Y�$��{� ���t�������p� �@���)�;� M���f�x����������� �����
.@@Rdv��,e� ����(: L^p�����`�� //��SK����!"�R/d/v/j�C]���  x/��/(� -$�����/z�)(���!O�*��C=pC?L?[��9  �?�65?�?�?�?��O �O9OKO]OoO�O(�U�O�O��O �O�O__'_9_K_]_ o_�_�_�_�_�_�_�_��_o#o/T1SV�GUNSPD�� �'u��F`2MO�DE_LIM �'��y�Bd2O`oa�(��AeASK_OPTIONj��y���a_DI��EN�B  ��u��aB�C2_GRP 2�)5%u�����@C��"s:lBCCFG' +�k(��2*�Yz`w����� ��	��-��Q�<� u�`�r�����Ϗ��� ޏ��'�M�8�q�\����������ݟ�$� ڜ	�۟<�N�ɟ+��� o�����̯ڪ5%�� ������>�,�b�P� ��t��������ο� �(��L�:�\ς�p� �ϔ��ϸ������� � �H�.��\�nߌߞ� ��.�������
���.� @�R� �v�d���� ����������<�*� `�N���r��������� ����&68J �n�Z߼��� �4"DjX� �������/ /./0/B/x/f/�/�/ �/�/�/�/�/??>? ,?b?P?�?t?�?�?�? �?�?O�O.OLO^O pO�?�O�O�O�O�O�O  __�O6_$_Z_H_~_ l_�_�_�_�_�_�_�_  ooDo2oTozoho�o �o�o�o�o�o�o�o
 @.dO|��� �N���*��N� `�r�@���������ޏ ̏����8�&�\�J� ��n�������ڟȟ�� �"��F�4�V�X�j� ����įzܯ��� 0���T�B�d���x��� ��ҿ�������>� ,�N�P�bϘφϼϪ� ��������:�(�^� L߂�pߦߔ߶߸���  ���$�گ<�N�l�~� ������������  �2� �V�D�z�h��� ������������
 @.dRt��� ����* `N�:���� �n//$/J/8/n/�X&� �$TBCS�G_GRP 2,�X%� � ��  
 ?�  �/�/�/�/�*�� ?">?E?/?�i?{=�"�#.�,d����1?�!	� HC� {6&�ff�2� {5�1A�x�!�?�9D)�{6���F|4AB4�?�?HL@YA�8$By�:O�MCj��PN�333{5B�C�O�O�O{9�O_��N|4>�G�AB�_Z]@�8[6�8�U�_ ^_p_�_�_�_�_o#o�2kh�La	V3�.002b	rc;2l2c	*n`fd��"}o<fG�?��33� X�ai 8�`�m�o  �# _X�o�e�!J2�#/�-��o
xCFG �1X%�!�!4z���"�b4�x����za �� ���+��O�:�s� ^�p�����͏���܏ � �%�K�6�o�Z��� ~�����۟Ɵ؟��� 5� �Y�k�q��v��� ��D�ͯ��ݯ��'� �K�6�o�������`� ɿ���ؿ��#ό!x/ H�T/X�Z�lϢϐ��� ����������D�2� h�Vߌ�z߰ߞ����� ��
���.��R�@�v� d���������� ��0���P�r�`��� ������������& 8��HJ\��� �����4" DFX�|��� ���
/0//T/B/ x/f/�/�/�/�/�/�/ �/??>?,?b?P?r? �?B��?�?�?~?O�? OO(O^OLO�OpO�O �O�O�O�O _�O$__ 4_Z_l_~_8_�_�_�_ �_�_�_�_ oo0o2o Dozoho�o�o�o�o�o �o�o
@.dR �v������ �*�<��?T�f�$�"� ����̏����ޏ �� �J�\�n�,�~����� ȟ������"�ܟF� 4�j�X�z�����į�� �֯�����0�f� T���x�����ҿ��� ���,��P�>�t�b� �φϘ���H�����
� ��:�(�J�p�^ߔ߂� �ߦ����� ����6� $�Z�H�j����n� ���������2� �V� D�f���z��������� ����
R@v d������� <*`rߊ �"�X��/�&/ /6/\/J/�/�/�/b/ t/�/�/�/�/"?4?F? X??|?j?�?�?�?�? �?�?�?OOBO0ORO xOfO�O�O�O�O�O�O �O�O_>_,_b_P_�_ t_�_�_�_�_�_o~ �.o@o�_o^opo�o �o�o�o�o�o$6 HlZ|~�� ���� ��D�2� h�V�x�z������ ԏ
���.��>�d�R� ��v�����П����� ��*��N�<�r�`��� ��Ro��ү䯎��� 8�&�H�J�\������� ȿڿ쿪����4�"ϜX�B�  ~���� �Ɩς��$T�BJOP_GRP� 22J��  ?���i	�µ�4���R�� �� ��,^�� ��� � s� � ��� �@~���	 �C�� 2�Qp�Dㄈ����N�&ff�V�K�W�i�<9]�2�?��?L��͊�BH  A�xHץ߰�D)���.>��SF�Y�����g��� �ҏ�>����<����?3�33?fh��B��  B ��=���D5mF��n�w�����Af������C+�&�.���Cj������߁����;ć�B��
�Ⴔ���]�����x�����<��6����F���j�|�NրO��"(����z��J6���>���C4(���}�� ������� &@*\f�r�������'/����ưJ!N�	V3�.00��rc2l��*t ��}��/��' F�  �F�  GX �G7� GR� �Gr0 G�� �G�@ G�� �G�\ G�� �G�` G�� �H
� Hd �H" H.� �H;� HH2 �HUޝ"E�� �E� �!F@ F�� Fj` F��� F� �"�!� G$ G� �GVص#�� G��L G�� G��h G�� =u=+,	XZ5���r?�2��=�3?�  &��~��ESTPAR �v�����HR�0A�BLE 15��# �0�0DD����|:�'�(P�(�ǉ��'	�(
�(Q�(A���(�(u�(�6RDI�?���FA����7OIO[OmH�DO�O�K�O_� _2_D^�2S�O��  �Joo)o;oMo_oqo �o�o�o�o�o�o�o %7I[���P�_ ��C�}�_�_�_�_gO�yO�O�O�O�H�2�rN�UM  J�*��"��� @�@��2_CFG 6�k��&�@��IMEBF_TT�1����0��VER�CAÆ���R 17Kg 8/�� ��fP�
 M��  � ��*�*�)�;�M�_�q� ��������˟ݟ�� �\�7�I���m���������ǯٯ���  �PDT�&� � "1[L�^� �{�M!������UK���ѿ�_�DE��� �OTF8,�>� �$Cd�v� �$�ϲ���s8�����RID��R�_e�چ@��0MI_CHAN��� � ��DBGL�VL����1��E�THERAD ?��5����00���:e��4:71:d0:66 ��m7��68�69��oROUT׀!iZ�!<�Z��9��SN�MASK������255.��2.�`#���5�����0O�OLOFS_DI� Tռ�ORQC?TRL 8��PS�?8�T'�\�n����� ������������" 4FXj|�K��؟��2PE)�TA�I����PGL_C�ONFIG >�k�{���/ce�ll/$CID$/grp1�M_q��KS���� ��//�>/P/b/ t/�/�/'/�/�/�/�/ ??�/�/L?^?p?�? �?�?5?�?�?�? OO $O�?HOZOlO~O�O�O 1OCO�O�O�O_ _2_�~}�Oh_z_�_�_�_ �_0���_�]��Oo 1oCoUogoyo�O�o�o �o�o�o�o�o-? Qcu���� ����)�;�M�_� q��������ˏݏ� ����7�I�[�m�� �� ���ǟٟ���� ��3�E�W�i�{����� .�ïկ������� A�S�e�w�����*����ѿ�����+�&��User V�iew ;}}1�234567890\�nπϒϤ϶Ͼ�XG�����B�2O� �� �2�D�V�h�z�����I�3��������� �"��C���4��|� ��������5�����5k�0�B�T�f�x��������6�����@,>��_��7�� ������Q��8�L^p����� l�Camera M�C//0/B/T/f/DRE��/�/�.Z��/��/�/??(?�   ���x?�?�?�?�? �?y/�?OOe?>OPO bOtO�O�O����� /O�O�O__,_>_�? b_t_�_�O�_�_�_�_ �_o�O�Gj�_Pobo to�o�o�oQ_�o�o�o =o(:L^po �GD;	����� ��o<�N�`������ ����̏ޏ����s� (�:�L�^�p���)��� ��ʟ�� ��$�6� H�G�	ߟ������ ʯܯ��$�6��� Z�l�~�������[��G :K� ��$�6�H�Z� �~ϐϢ�������� ��� �ǿٷ9��a� s߅ߗߩ߻�b����� ���9�K�]�o����"	�0����� ����(���L�^�p� �������������� ������GYk} ��H����4 1CUg�[; ������/� 1/C/U/�y/�/�/�/ �/�/z���Kj/?1? C?U?g?y? /�?�?�? ?�?�?	OO-O?O�/ �%3k�?�O�O�O�O�O �O�?	__-_xOQ_c_ u_�_�_�_RO�%�{B_ �_	oo-o?oQo�Ouo �o�o�_�o�o�o�o �_�%��ocu� ���do���P�)�;�M�_�q���*}  .y��ď֏� ����0�B�T�f�x��   � b��Ë!��L���?�-A�
��C�b*qDlN�Ø@P�y���@6��@��ߦ�1�∍?�łBl@֑v������z�ǟ Aǒ^�"�\�D�H�ɿ
D;��Ғ??u�C%R,Z��� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϰ����������*p
*p(  �覀( 	  ��0��T�B�x�fߜ� �߬߮���������t>�,��� �� ������������ �%�,sr�O�a�s��� ������������8� '9��]o��� ������F#5 GYk}���� ��//1/C/U/ �y/�/�/��/�/�/ �/	??b/??Q?c?�/ �?�?�?�?�?�?(?:? O)O;O�?_OqO�O�O �O�O O�O�O_HO%_ 7_I_[_m__�O�_�_ �__�_�_o!o3oEo �_�_{o�o�o�_�o�o �o�odoASe �o������* ��+�rO�a�s��� ������ߏ��J� '�9�K�]�o���ȏ�� ��ɟ�����#�5� G���k�}���֟��ů�ׯ����T�4�@ A/�<�N�`�/�6�����)frh:�\tpgl\ro�bots\r20�00ic��_12?5l.xml�Ŀ ֿ�����0�B�T�f�r���rϗϩϻ� ��������'�9�K� ]�t�nߓߥ߷����� �����#�5�G�Y�p� j������������ ��1�C�U�l�f��� ������������	 -?Qh�b��� ����); Md^����� ��//%/7/I/` Z//�/�/�/�/�/�/��/?!?3?E?W>y�ί� 6���<<w �� ?�W; �?W?�?�?�?�?�?O �?0ONO4OFOhO�O|O �O�O�O�O_�O�O_�J_X��$TPG�L_OUTPUT� Ab�b�� z0C��b��2�D����?�-B^}��C6�q^�ê�Dó B^�@6���B��P1�� ^��_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7Ewz0��OPcell/c�ont1/grp�1/dcs/cp�cz/z6/f ��eB��� ��,kB�PX��q� ��g�R����X�7�@^����� �QBУ��X��u^��p�CXO�r�u[mx1y�u��p�q�ZOB�X��$A�R�u���֊s<���v23�45678901 f�x���������ȃ�s d�����&�8�J��s}M�u���������U� g����)�;�M�� [���������˯c�ٯ ��%�7�I���� ������ǿٿq��� !�3�E�W��eύϟ� ������m����/� A�S�e���sߛ߭߿� ����{����+�=�O� a����������� �����'�9�K�]�o�׍}u1�������������
@|?.@�:? ( 	 Cu c������� �;)_M�q �����/�%/ /I/7/Y/[/m/�/�/�/Qv�x0�6�/?= �/5?G?!?k?}?Kz�/ �?�?Z?�?�?�?�?,O >O�?BOtOO`O�O�O �O�O�OPO�O(_�O_ ^_p_J_�_�__�_�_ �_�_o$o�_0oZo�_ �_�o�o<o�o�o�o�o  ~oDV�oB� fx��2�
�� �@�R�,�v����p� ��Џj������<� ��$�r���������� ���N�`�&�8�ҟD� n�H�Z��������� ��د"�4��X�j�ȯ R���:���ֿ�¿� �|��T�f� ϊϜ� vϨ���0�B��ߴ� "�P�*�<߆ߘ��ϼ� ��hߺ������:�L���")WGL1.�XML
���$T�POFF_LIM� �  �!����N_SV�� � ��P_M�ON B�%ԫ�  2��ST�RTCHK C��%������VTCOMPAT��H���VWVAR Dr��k��� �� �� ����_�DEFPROG �%�%PN�S0001 IO?NCHECK�����_DISPLAY������INST_�MSK   ���INUSER�>���LCKGQUICKMENk���SCRE� ��%I�tpsc@��G� �	�� _�	�ST<���RACE_CFG E���k���	��
?��HNL 2F��� *r� ��^p �������ITEM 2GJ� �%$12345678901/C%  =<;/a/s/{#  !�/�+��E/�/��//�/S/? %?�/;?�/�/�?�/�? ?�?�?_?O?a?s?�? �?O�?gO�O�OO�O 'O9OKO�OoO_A_S_ �O__�O�O�O�_�_5_ �_ok_o�_�_jo�_ �o�_�o�oo�oCo�o yo9�oIo��o �	-�Q�#� 5��Y����e�}� �׏�M���q���L� ��g�ˏ�������%� 7� �[���+�Q�ן ǟٟ�����3�߯ ��{�;�����ï=� 篓���˿/�׿S�e� w���Iϭ�m��㿋� ����=���a�!�3� ��I߻�ߖ��ϱ�� ������]��ߓߥ� ���u������5� G�Y������O�a��� m����������C��y�+����xS�H}
�  �}
 "���
 ��+�
�UD1:\8����R_GRP �1I+� 	 @_ ��� ������ $/�2*�8\/G/�/k%?�  �/�+�/�/�/ �/�/??%?'?9?o? ]?�?�?�?�?�?�?�?�O	K%O7O�S�CB 2J� �/�O�O�O�O�O�O��O__�UTOR?IAL K��^_�V_CONFIG L�z��_n\OUTP�UT M�	�P���_oo1oCo Uogoyo�o�o�o�o�o��o_�\Reg�ular Option�o0BT fx����������_�!�3�E�W� i�{�������ÏՏ� �d��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v������� ��п����*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x�����������������U� ���_9K]o�� ������� 5GYk}��� ����/1/C/ U/g/y/�/�/�/�/�/ �/�/	??,/??Q?c? u?�?�?�?�?�?�?�? OO(?;OMO_OqO�O �O�O�O�O�O�O__ $O7_I_[_m__�_�_ �_�_�_�_�_o!o2_ EoWoio{o�o�o�o�o �o�o�o.oAS ew������ ���*=�O�a�s� ��������͏ߏ�� �'�8�K�]�o����� ����ɟ۟����#��C�B�J�X��>�-��"\Re�gular Option����ί� ���(�:�L�^�p� ��5�������ѿ��� ��+�=�O�a�sυ� 6��ϻ��������� '�9�K�]�o߁ߒϥ� �����������#�5� G�Y�k�}��߳��� ��������1�C�U� g�y������������ ��	-?Qcu �������� );M_q�� �����//%/ 7/I/[/m//�/��/ �/�/�/�/?!?3?E? W?i?{?�?�/�?�?�? �?�?OO/OAOSOeO�wO�O�O�$TX_�SCREEN 1}NV�>��}��O�O�O__(_:_�O���Oz_�_ �_�_�_�_K_]_
oo .o@oRodo�_�o�_�o �o�o�o�o}o*�o N`r���1 ����&�8��\� ���������ȏڏQ� ��u�"�4�F�X�j�|� ����ğ֟���� ��0���T�f�x��������%�ү�$UAL�RM_MSG ?5�I��@ ʯ�: ��G�:�k�^����� �������ܿ� �1�~�SEV  ��c��ECFG� P�E�A � �5@�  A���   Bȧ1�H�@�����l� �A �XT�e����TɈ3~����Tɖ\�Ͽ�gT�S�����T�$�
�!	�qT�am
��5�T�e�:���T��u�R���T���j��T�B��o�GRP 2Q�y� 0��	 �����k���
����"���x|������:�I_BBL_NOTE Ry��T��lȧ2�@�1����DE�FPRO�%�� (%PLAC�E_<�STIC_�PALLET_L�EFT�:%CL?EAR_IO2�V� %Ϝ�������������,�>�)�b���FK�EYDATA 1�S�I  	p 9�ǟ6 h���`��������,(�=�4+ OINT�]�EG OOK T����tNDIRE�CT��TCHOI�CE`�X UCH�UP��X RE INFk�#`rY �}�����/�&//J/1/n/�/�����/frh/g�ui/white�home.png��/�/�/�/�/?� } �%point�/�<?N?`?r?�??/look+2.1.?�?�?��?�?O8indirec*?FOXOjO|O|�O>choic�#if�O�O�O�O__�8touchup�6ON_`_r_�_�_>arwrg5O�_�_�_ oo�X5oGoYoko}o �o�o0o�o�o�o�o �oCUgy�� ,����	��-� �Q�c�u�������:� Ϗ����)���M� _�q����������%�� ���	��-�?�F�c� u���������L��� ��)�;�ʯM�q��� ������˿Z���� %�7�I�ؿm�ϑϣ� ����V������!�3� E�W���{ߍߟ߱��� ��d�����/�A�S� ��e��������� r���+�=�O�a��� ������������n��� '9K]o���@������+��� �4F�""o��#,g/�_(OPY   ]�~� OOK L��/�AD D T�// AVE A�S9/:/  RINT Pe/f/�/�/�/ �/�/�/?�/3??W? i?P?�?t?�?�?�?�?�Ɲ&Ewhitehom�CO1OCOUOgO<v,Wpoin�_�O�O�O�O�O�Oi/look�B�O4_F_X_�j_|_�Lindirec�O�_�_�_�_�_>�NchoicC�_�>oPoboto�o�Jtouchup�_�o�o��o�o�Narwrg�_@Rdv� �������*� <�N�`�r�����%��� ̏ޏ������8�J� \�n�����!���ȟڟ ����"���F�X�j� |�����/�į֯��� ���?��T�f�x��� ������ҿ����� ,ϻ�P�b�tφϘϪ� ��K�������(�:� ��^�p߂ߔߦ߸�G� ���� ��$�6�H��� l�~������U��� ��� �2�D���h�z� ����������c���
 .@R��v�� ���_�* <N`����� ��m//&/8/J/�\/3�j+�@ j/�/�/B�/�/�/ C�,�??�8OINT�  ]%?'? IR�ECT Q?R?  �NDf2}?? CH�OICE@?�?80UCHUP�?�?O%O OIO0OmOOfO�O�O �O�O�O�O�O!_3__�W_6��Uwhitehom'c�_�_�_�_x�_�gpoin/�o-o?oQoco�_i/direc
o�o�op�o�o�owo/in�o�!3EWi�oachoic�_������/touchup�.�@�R�d�|v��^arwrg ��ԏ�����.� @�R�d�v�������� П������*�<�N� `�r��������̯ޯ ����&�8�J�\�n� ����!���ȿڿ��� ϟ�4�F�X�j�|ώ� e_+����������� %�B�T�f�xߊߜ�+� ����������,�� P�b�t����9��� ������(���L�^� p���������G�����  $6��Zl~ ���C���  2D�hz�� ��Q��
//./ @/�d/v/�/�/�/�/ �/_/�/??*?<?N? �/r?�?�?�?�?�?����;�sP���OO'M�?IO[O5F,G_�O?_�O�O�O �O�O
_�O._@_'_d_ K_�_�_�_�_�_�_�_ �_o�_<o#o`oroYo �o}o�o�o���o &8JY?n��� ���i��"�4� F�X��|�������ď ֏e�����0�B�T� f�����������ҟ� s���,�>�P�b�� ��������ί�򯁯 �(�:�L�^�p����� ����ʿܿ�}��$� 6�H�Z�l�~�Ϣϴ� �������ϋ� �2�D� V�h�z�	ߞ߰����� ����
��o.�@�R�d� v��߬�������� ����<�N�`�r��� ��%��������� ��8J\n��� 3����"� FXj|��/� ���//0/�T/ f/x/�/�/�/=/�/�/ �/??,?�/P?b?t? �?�?�?�?K?�?�?O O(O:O�?^OpO�O�O �O�OGO�O�O __$_h6_H_�J[�����s_�_�]o_�_�_�V,�o�_�o  ooDoVo=ozoao�o �o�o�o�o�o
�o. RdK�o�� �����*�<�� `�r����������Oޏ ����&�8�J�ُn� ��������ȟW���� �"�4�F�՟j�|��� ����į֯e����� 0�B�T��x������� ��ҿa�����,�>� P�b��ϘϪϼ��� ��o���(�:�L�^� �ςߔߦ߸������� }��$�6�H�Z�l��� ����������y��  �2�D�V�h�z�Q��� ������������. @Rdv��� ����*<N `r����� �//�8/J/\/n/ �/�/!/�/�/�/�/�/ ?�/4?F?X?j?|?�? �?/?�?�?�?�?OO �?BOTOfOxO�O�O+O �O�O�O�O__,_�O P_b_t_�_�_�_9_�_ �_�_oo(o�_Lo^o@po�o�o�o�o���k���������o�o}�o);v, '�l��w��� ��� ��D�+�h� z�a�����ԏ���� ߏ��@�R�9�v�]� ������П����� *�9oN�`�r������� ��I�ޯ���&�8� ǯ\�n���������E� ڿ����"�4�F�տ j�|ώϠϲ���S��� ����0�B���f�x� �ߜ߮�����a���� �,�>�P���t��� �����]�����(� :�L�^���������� ����k� $6H Z��~����� ��� 2DVh o������� �/./@/R/d/v// �/�/�/�/�/�/�/? *?<?N?`?r?�??�? �?�?�?�?O�?&O8O JO\OnO�OO�O�O�O �O�O�O_�O4_F_X_ j_|_�__�_�_�_�_ �_o�_0oBoTofoxo �o�o+o�o�o�o�o �o>Pbt�� '������(��� *��� ���S�e�w�O�������,��܏�� �� $�6��Z�A�~���w� ����؟�џ���2� D�+�h�O���s���¯ ���ͯ
���@�R� d�v��������п� ����*Ϲ�N�`�r� �ϖϨ�7�������� �&ߵ�J�\�n߀ߒ� �߶�E��������"� 4���X�j�|���� A���������0�B� ��f�x���������O� ����,>��b t�����]� (:L�p� ����Y� // $/6/H/Z/1�~/�/�/ �/�/�/��/? ?2? D?V?h?�/�?�?�?�? �?�?u?
OO.O@ORO dO�?�O�O�O�O�O�O �O�O_*_<_N_`_r_ _�_�_�_�_�_�__ o&o8oJo\ono�oo �o�o�o�o�o�o�o" 4FXj|�� ������0�B� T�f�x��������ҏ ������,�>�P�b��t�����o ���>o ���ß՟ 睿�	����,�L� ��p�W�������ʯ�� � ��$��H�Z�A� ~�e�������ؿ���� � �2��V�=�zό� k/����������
�� .�@�R�d�v߈ߚ�)� �����������<� N�`�r���%���� ������&���J�\� n�������3������� ��"��FXj| ���A��� 0�Tfx�� �=���//,/ >/�b/t/�/�/�/�/ K/�/�/??(?:?�/ ^?p?�?�?�?�?�?�� �? OO$O6OHOO?lO ~O�O�O�O�O�OgO�O _ _2_D_V_�Oz_�_ �_�_�_�_c_�_
oo .o@oRodo�_�o�o�o �o�o�oqo*< N`�o����� ���&�8�J�\� n��������ȏڏ� {��"�4�F�X�j�|� �����ğ֟����� �0�B�T�f�x���������ү�����0�
���0���3�E�W�/�y���e�,wϼ�o��ǿ�� ��:�!�^�p�Wϔ�{� ���ϱ������$�� H�/�l�Sߐߢ߉��� �������? �2�D�V� h�z��������� ��
���.�@�R�d�v� ������������� ��*<N`r�� %����� 8J\n��!� ����/"/�F/ X/j/|/�/�///�/�/ �/�/??�/B?T?f? x?�?�?�?=?�?�?�? OO,O�?PObOtO�O �O�O9O�O�O�O__ (_:_�^_p_�_�_�_ �_�O�_�_ oo$o6o Ho�_lo~o�o�o�o�o Uo�o�o 2D�o hz�����c �
��.�@�R��v� ��������Џ_��� �*�<�N�`���� ����̟ޟm���&� 8�J�\�럀������� ȯگ�{��"�4�F� X�j���������Ŀֿ �w���0�B�T�f��x��$UI_IN�USER  ��������  y�}�_�MENHIST �1T�� � ( �����'/SOFTP�ART/GENL�INK?curr�ent=menu�page,74,�1 1 TE�VERIFY�)�;��M�_��)���16�31�ALLET_LEFT�ШҐ��������(v߈�4�8,2  ,59� ��HEIGHT?_CHECK��I��[������7�� P�LASTIC_P���9������߁��8���PROGRAM �/�H�Z�l�w����34,4 _JACKPO�ѡ�@�=������s�4����ed�it�JR_SETU,����Ugy<t�,HOMѰ�p;���� ��� ��.@Rdv� ����� /�+/=/O/a/s/�/ /�/�/�/�/�/?? �/9?K?]?o?�?�?"? �?�?�?�?�?O�?5O GOYOkO}O�O�O0O�O �O�O�O__
C_U_ g_y_�_�_�_�O�_�_ �_	oo-o�_Qocouo �o�o�o:o�o�o�o );�o_q�� ��H����%� 7��[�m�������� ǏV�����!�3�E� 0_N�{�������ß՟ ؏����/�A�S�� w���������ѯ`�� ��+�=�O�a�𯅿 ������Ϳ߿n��� '�9�K�]��nϓϥ� ��������|��#�5� G�Y�k�V�ߡ߳��� ���������1�C�U� g�y���������� ��	���-�?�Q�c�u� ������������� ��);M_q�� $������7I[m�|���$UI_PANE�DATA 1V������  	�}c/�frh/cgtp�/flexdev�.stm?_wi�dth=0&_h�eight=10���ice=TP�&_lines=�15&_colu�mns=4�fo�nt=24&_p�age=whol�e��z�)prsimA/j/  }m/��/�/�/�/�/�/ ) �/?�/5??Y?k?R? �?v?�?�?�?�?�?O�OOCOz����    %"Ҷ{$����2
%3�@.1(%d�oub�@2MO+Hu�al�O
_qKitree�A_E_W_i_{_ �O�_�_�_�_�_�_o �_/ooSoeoLo�opo��o�o�o�oVH bC? m�X�sO�O�OP3
&( �O(%�t#p3�o�khird��~/���� �)��oM�4�q���j� ����ˏ��ݏ��%���I�[�B���odA? 	2W�.t�� ǟٟ����b�!�E� �i�{�������ï*� �ί����A�(�e� w�^�������ѿ����ܿ�+��bB��_� d�vψϚϬϾ���� U���*�<�N�`��� �ߖ�}ߺߡ������� ���8��\�n�U�� y����;�M����"� 4�F�X���|��Ϡ��� ��������s�0 T;x�q��� ���,>%b ��������� E/(/��L/^/p/�/ �/�//�/�/�/ ?�/ $??H?Z?A?~?e?�? �?�?�?�?�?o�?/ DOVOhOzO�O�O�?�O 5/�O�O
__._@_�O d_v_]_�_�_�_�_�_ �_�_o�_<oNo5oro Yo�o�oO-D��o�o �o
.@)�oe �ET������ R��3��,�i�P� ��t���Ï���Ώ����A��H+C%K�$�UI_POSTY�PE  +E�� 	 ��`�� �����Cs�Q�UICKMEN ; �� �����_RESTOREw 1W+E����*de�fault�K � OUBLE��PRIM�m�editpage�,JR_SETU�PPROGRAM�,1N�������T�omenuf�98z� � ��$�W�.�R�d� v�����-�4�����/� �
��.�@�R���v� �ϚϬϾ�a������ �*�տ7�I�[��ϖ� �ߺ����߁���&� 8�J�\��߀���� ��s�������k�4�F� X�j�|���������� ����0BT�� 	s������� �>Pbt��)�������S�CRE?ǝ�u1sc��u23$33$43$5*3$63$73$83!#wTAT~�� ֓<+Ek�USER /�,$ks5#�$3�$4��$5�$6�$7�$8��!s�NDO_CFOG X����s��PDv!�)��None��� _INFO 1Y+E5Z0Ԑ0%�u? �Hc?�?�?�?�?�?�? O�?4OOXOjOMO�O�O�O�O��G1OFFNn� \��^1�O ���_'_9_K_x_ o_�_�_�_�__�_o �_o>o5oGotoko}o@�o�[ן�m�o�o
�oL#�HUFw�7���6D1RTOL_�ABRTGB3_rE�NBhYxGRP �1]�ӑCz  A��s�q1�� ����(�:�[v���U�x1w{MSK � �uZ1���[vN�Dq%R9�%P�NS000ޯ.RO_EVNgp��6��22^�K
 h�1UEVgp!�td:\eve�nt_user\�Џ+�C70� 0F�e�#�SP)�.�spotweld`�!C6��f�x���d!�o?���2�ݗ�� �!��e���E�W�Я {�������ï<��`� ��S�����̿w��� ����8����n�� �Ϥ�O�a��υ��ϩ���� �WRK 2_��)q8��b�t�  Pߙ߫߆����߼�� ���;�M�(�q��^� �����������%�� �6�[�m��$VA�RS_CONFI�0`�K FP���t�CCRG2�c�J�O����D,A��BHJ�p�C�J��*(?��: �$��MR�r2iN�Kl�0	q����@1: SC�130EF2 *(�� ���X��ș�˂501<A@vC��� ���!Ns�Iv�8�,0�b� B�����Z�: /�;/&/_/J/�/n/ �/�//�/�/�/�/%?p�I?[?��TCC��j�z@�98���j ���GF��
�k�K� �%UF12� Auto �0 �e set ��R� �h?"u 
�1�em�~3456?789012I��A� �0������H�������fX:���3��.:$@8�@�9� (:�o=L�m���y����%I��O��j����%���O��1 ��_%W[B-hOzO�O �O�_�O�H�_�__%_ '_9_K_]_o_�_no�_ �_�o�_�_�oo#o5o�Go~�1SELEC�넙����qVIA�_WO:�l��|�p��,		��`|�o�G�P ǫp��iXqSIONTM;OU� ��u���m�:��<�t�1 FR:}\�s\DATA̟��0�� UD1w:\ �LOG��   %��EX�0�' B@� ��s�D�  �1.200.��5�2 .design.local;��[���= �� � �n6  ���8��p��t#`φ	  =�������� 
 MC>�vTRAINZ��24��dO�p�����m�}��sOn�; (1[���
9���� ��џ���=�+�E��O�a�s�����z�ISSTAT o�9�y� =-2997�.6665: w�as less �than acc�eptable �value: -�1��0)���$80_?SIDE_B4�g;_IS_GE�sp�;����
rpj ���\�HOMIN�pq/�E�����rq$q�aC$B�m\��JMPERR 2=r�;
  �o�� ���e���.�_�R�d� vψϚϬ�������ϰ�Dc�W�RE�ps\�|�LEXg�t����@1-eP�VMPHASE  ���j!r�OFFS_ET_ENB��u�OyP2�tu�F%��|���<cB�`A�1�`� ?s33���1cA��cEP��|��x��H��x��A �t�^ �= ��b�3������I�?��i� �����Õ������3�,�?5�����r� �օ�&��Z��w?� 1����Ⱦ��{�1��� ����!S���#��~ �������+  OAsh��� ����
/9K ]R/�'/�/�/�/ �/�]/�/5/*?<?k/ ]?�/i?�?�?�/�?�/ �??OC?U?�?EOSO eO{O�?�O�?�?	O�O -O�O�O+_=_O_y_�O 	_{_�O�_�__	os_ o?o9o�_xo�_�o�_ �o�_oKo�o�o'�5w[�TD_FIL�TE�yo� �g�t����o��� �����'�9�� �f�x���������ҏ�����W�SHIF�TMENU 1z�<�%�f�1� D�j���z���ٟ�� �����W�.�@����d�v�ï��	LIVE/SNAP��vsfliv���կ�b�ION� ��U���menu����r���3�$�j��{b���MO���|n��zY�WAI�TDINEND � ��Kᷲ�OK�����OUT��S�,���TIML���W�G�y�Ϝ�+��|�J�|�i���REL1E������TM�˳�{��_ACT����u���_DATA� }b�v�%  �RIPPER_O�PEN���`�RD�IS1�-��$X5S��~b�����J���Z�XVR���;�$ZABC_GRP 1��ٕ�`,�h2���ZIP���F�sc�o������z�MPCF�_G 1��� A0�o'���?�����`p�� 	|�y�  <T��  7�?���;�Tؿ���7�{�����ֺ������T���D�^�@C2�{q�0f������jD� �����x�������  4��A��Sa���7Q�v��������SF������?�qC2��wa����k���
����"���|����?���k^|�f���b �����򘾹ϝ-B��!��?޿�������o ��
 .X�������cN��������� I�" p�& �:.�>,�w��ৰ����_C_YLINDfq���� Јf ,(  */.-�c/W/>/{/b- ��/�/ �./�/g/???R? �/v?�?�?�/�?Y??? �?�?O�?m?NO`O��?�2���x� � ��O�o��O�_\h�O8_�g�RQA���SPHERE 2��̲?�_O�_�_ �_�_0OC_o0o�?To �_�_�oqo�o�oo�o �o=oOo,�oP7I���o���9�ZZ�� ǳ�