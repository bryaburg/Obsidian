��   �A��*SYST�EM*��V9.1�0170 9/�18/2019 A 	  ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTTR_&F/�� $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STSTOP�_TPCHG �V LOG_P NT��N�  6 C�OUNT_DOW�N�$ENB_�PCMPWD� �$DV_� IN�� $C� CR5E��A RM9� =T9DIAG9(|�LVCHK >FULLM/��YXT�CNTD��MENU�A�UTO+�FG_wDSP�RLS��U�BURYBA�N�!  &EN}C/  �CRYPTE ����$$CL�(   ����K!�� T @ V� I�ONH(; ��Z�$DCS_7COD?���O%��H ^z'_� �-]W�(S  J*�� IL �&�A91�"�K!	 
 $R!��=?$? 2?H?V?l?z?�?�?�? �?�?�?�?
O O.ODO\<#'SUP� �*a�FOXO�#FxO��O�O��  ��L�A��_ � ��� V�[t&�+�j���D�O`_ ��W_��;!�U�_cGLUGH 1K)_ ; �) �_�_	oo-o?oQoco uo�o�o�o�o�'�_�o �o!3EWi{ �����o��� �/�A�S�e�w����� ����������+� =�O�a�s��������� ͟܏���'�9�K� ]�o���������ɯ؟ د���#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ��������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi{ �������%