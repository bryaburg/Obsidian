��   ��A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����DCSS_C�PC_T  �4 $COMM�ENT $�ENABLE � $MODJG�RP_NUMKL�\  $U�FRM\] _VT�X M �   �$Y�Z1K �$Z2�STOP�_TYPKDSB�IO�IDXKE�NBL_CALM�D�USE_PR�EDIC? �EL�AY_TIMJS�PEED_CTR�LKOVR_LI�M? p D� L�0��UTOOi��O�  &S. ǰ 8J\TC �u
!���\�� jY0 � � �CHG�_SIZ�$A�P!�E�DIS"�]$!�C_+{#�s%O#J�p 	]$J d#� �&s"�"{#�)�$��'�_SEEX�PAN#N��,$STAT/ �DFP_BAS�E $0Kf$4!� .6_V7>]H73��&J- � }�\7AXS\UP��LW�7����s�$d4r �<  w?�?�?��?�?�/x/) jELEM/ T �&B.2�NO�G]@%CNHA��DF#� $DAT�A)he0  �PJ�@ 2� 
&P5 �� 1U*n   �_VSiSZbRj0jR(��VyT(�R%S{TR/OBOT�X�SAR�o�U�V$CUR�_��RjSETU�4"	 �bAISP�_MGN�INP_ASSe#�PB! � `CiH�77`e�.f�Xc1�CONFI�G_CHK`E_P�O* }dSHRST�gM^#/eOTHEoRRBT�j_G]�R�dTv �ku�chT1r
0R HLH�d� 0  lt<Ne'AVRFYhH^t�5"�1� ��W�_A�$R�4SPH/ (G%Q��Q�Q3wBOX/ 8�@F!�F!��G �r{�sc4TU�IRi@  ,��F�pER%@2� $�p �L�_SF��eUI�ZN/ 0 �IF(@�p��Z_��0�_�0wu0 � @�Q7yv	
��~ � �$$CL` � ��a0�����Q��Q��VER�SION���  �Z�$�' 2 �Q � Cel�l Box In8��*�h� ���m����PE"�� œ�����E�� ŷ�����ĨO� D�ğ�����  d����Cz � ����:���JackpotT�Out_�q�w�������c��@����^π DH��Κ�@�ȯ+���9�'�I��Incoming�[�n�����a  E�	����D\  �ȩ���ޡ�ÿ-�� �;�)�G�H�l�{��� oϬ�������h����%�7�I�Midd�leT�h�~���9 � �8`L߫�C��&få��Οl�
��	2���@�>�D��Left Si�de�`�u��ߐ�;� E�߭�CԐ����>Д�  D����с����D�B�D�Righg�z��� �����ྱ������Q���%�K�9O�IC�K SLOWDO�W�z�߃�ؐ��������ě�����n�0BWb��d�J2 SlowdowZ�������&�����[�Cې�����1/E/_��h�z����D �����/#/5/ ?I?Sπ?wωϿ��? �?�?�??1?C?U? g?|O�O�?�?�O�?�O �O�OO-O?OQOf_Y��pick dcs tesb��)����_��Ö@P�P�_`��ې�Qo_._@_ R_TorO�o�O�O�O�o �o�o	o*o<oNo`o ro���o�o��o� ��&8J\�� ����p��̏�� "�4�F�l�j�|���� ��ďٟ�����0� B�T�f�{��������� ������,�>�P� v�d���������ί� ���(�:�L�^�p� �ϔ��ϸ�ʿ���� �'�6�H�Z� �nߐ� �ߴ����������#� 2�D�V�h�zߏ�߳� ����������1�@� R�d�v�x�������� �����-<�N�`� r������������ )�J\n� ;������� %/7/FXj��� �/@/���//!?3? B/T/f/x/�/�?�/�? �/�/�??	O/OAOP? b?t?�?�O�?�O�?�? �?_O+_=_LO^OpO �O�O�_�O�_�O�Oo _'o9oKoZ_l_~_$o �o�_�o�_�_�_ o 5GVohozo�o�o� �o��o�o�1�C� U�dv�����ӏ ��*��
�?�Q�`��r����������$D�CSS_CSC �2��ۑ�Q  P�100% Saf?e Spee}�b�.l�F@
,�ł{�j�d1��j�C���'�,�
����i�����d�����ԯ5��� Y��i���R���v�׿ ��������1�U�� y�<ϝ�`��τ����� �����?��c�&߇� J�\߽߀��ߤ���� )���9�_�"��F���j����ΔGRP �2ۛ �Ä�C��\Enњ�C  E5�� 	��5�ǀ#�\�G� ��k������������� ��F1jU� y������ 0T?xc�� ����/�/>/ )/b/M/�/�/�/u/�/ �/�/�/?(??L?7? p?�?�?_?�?�?�?�?  O�?�?6O!OZOlO~O IO�O�O�O�O�O�O_  __D_V_h_3_�_w_ �_�_�_�_�_�_�_.o�ŝGSTAT 2�ۙ-��<� ��?]����� 9�EL������]�����2F;��;���f��2D��J�O��DI�ۑ`<jf��;����Ɓ2%�=g4�t?��  �a��`4���ZC��@���Ɓۑje���S�<��?t�M��tg�<�ﾗ���i�Ʉ�@>F �D�Y�x�i>G[����0?}�}<����a��Ϳ�}��<���>�W�A�,]�9v�D�9]{�F�+�S?}۷)BsÊJq� �����.����D�.�U�zD~ܫ�i?�����;�~�=p�p.;�ϵ������˙?�b�no�o �o�gە�0�ە�\� n�H��������j�`i ҏk�z����	�+� -�?�a���u���ş�� ��ߟះ�=�O���[� ��_�q���ͯÏ��� %��-��%�G�u�[� }��������ǿٿ�� )�+�ѯkϝ�Wϡϳ����������?]�`��  �9�q��pq�]������;�X7;�뒌�p1�`�O�γDI��o��3��"�b2%TE��`�bS��`3�d�;�	+�o��<�#�`W�`�<�߸pNf���t >F@p�~{J��u>2p]<�"N�>p�6Bp�<��>�[YA�6���9��Vp_{ٯ�+��np	���G�ѽ"�p&�ϧ��p�U�&dD~�)�|���'C;}���=�p&;Ϫ5���Vٻː. �p1�(�
��.��Ϻ� �����������8�J� �2�t�Fό������� ��������(@^ DVx�L���� �0
Tf\�� �������/ �/D/*/</^/�/r/ �/�/�/n?6�/:? L?&?p?�?\?z��2� D�V�h�zߌߞ߰��� ������
��.�@�R� �O�?�?�?d?V_h_^? t_�_x_�_�_�_��/ o�/(oFo,o>o`o�o to�o�o�o�o�o�o�o B�/r��_p� �����_F,�Z $�F�t�Z�|������� ��Ə؏��(��0�^� D�
������֟� ����_(_�?�?�? OO(O:OLO^OpO�O �O�O�O�O�O�O`�B� T�f� ������:� �&�pς��j���~� ����������*��2� `�F�xߖ�|ߎ߰��� ��� �R��V�h�B� �������������� ����F�,�N�|�b� t��������������� <n�(r�^�� ���Ŀj�|������� į֯�����0�B� T�f�x������ ��/�/��/�/�/�/ ??��H?`?~? d?v?�?�?�?�?�?�? O2OO*OLOzO �O �O�/�O�O_�O(_:_ 0?~Od_�O\_~_�_�_ �_�_�_�_o�_o2o `oFoho�o|oB_�o
_ �o �oDV0N/ `/*<N`r �������/ /&/��z��8*� <�2H�r�L�^����� T_�o䟶o��� �� 4�b�H�j���~���ί ��Ư���oF�X��� D�����z�Ŀֿ̟�  �.����H�.�P�~� dφϴϚϬ������� �2��޿tߦ�`ߪ� �ߖ����������� ������ �2� D�V�h�z������� 4��(�:��������� ������DV�>� �Rߘ����� �4LjPb ��X���&�*/ <//`/r/h��/� �/�/�/�/�/? ?"? P?6?H?j?�?~?�?�? �?z/OB/�?FOXO2O |O�OhO����>�P�b� t����������� ��(�:�L�^��_�O �O�OpObotojO�o�o �o�o�o�o�/�?�? 4R8Jl��� ������ �N� �?~����o|�Ə؏�� ���R�8�f�0�R� ��f����������ҟ ��4��<�j�P�� ��ޏ�����ί�*��8��$DCSS_�JPC 2"��Q ( D�Right �Side Cle�ar����C9 W @@��
#P"QLefn��������Õ������In j�������C�*�� �����򰮶����!��/�"�`{�B�Ȏ��At Pick|���A  ����$�
RH Jac�kpot��̕�CD!���L�߇��a��ݳkό�Sߡ��Ⱦ�H?ome J1�����ٙ���ff�4���2�����O��������3����������3_�G���4a��%��������5���¤  ¤��r��6�����>����at E�OAT chg ����B�ffB��R�f��/�@Fff@����_�s�?���������8���&` ?�vߨ�t����b j��d���+�?�B�  B��bdsblB�� f����� �������2������$.�3J�
�'�"{4���"Q�����5 a��� �j��6��� �B�>/�ߥ/�߮�~F�2 limiO�V.�B�
�P���# ��/�/?#P�/m? �/�?`?�?�?�?�?�? �?�?3OOAO&O{OJO �OnO�O�O�O�O_�O �OA__"_4_�_X_�_�|_�_�_�_J�SS��W�L  afe? Speed�_»Bȉ�H�1aG�a2&`to�o7�A8�� aaai��ro�o�_�ofa �o�o?c*� N�r����� �;�M��q�8���\� ����ݏ���ȏ%�� 3��m�4�F�X�j�ǟ ��럲��֟3���W� �{�B���f�x���� ������A��e�,� ��P���t�ѿ��߿�� �����s�:ϗ� ^ϻς��Ϧ����'� ��K��$�6ߓߥ�l� �ߐ��ߴ����5��� Y� �}�D��h���� ��������C�
�g� .���R���v������� ������?Qu< �`����� )�7q8J\�n����dMO�DEL 2k�x^!��$<��c�X B���fÈ  A`�  CHp �� ��o$F/X/�	p xp$6  ë$�/�/j&�t(� �/�/�&�!�%�#�9�!�hM7 b?9?K?�?o?�?�?�? �?�?O�?�?LO#O5O<GO�WJ3 �O=-M=C\�(s �s 3��� �@CW�CbO tO�O\O__e_<_N_ �_r_�_�_�_�_�_o �_oOo&o8oWo\ono`�o�o�o�o� �L�o�o\�oEWi {������� ��/�A���e�w�ď ������я���B�� +�x�%S�e�ҟM� ��͟���P�'�9� ��]�o���ί����� ۯ�:��#�5���Y� k������������ ۿ�ÿ1�Cϐ�g�y� �ϝϯ���������D� �-�z�Q�c�u߇ߙ� ��������.���)� ����#�Q�c�9��� �����<��%�7�I� [�m������������� ����!nEW� {��u������ F/|Se�� �����0/// f/=/O/a/�/�/�/�/ �/�/?�/??�t? =?O?�?�?�?�?�? �?�?�?O#OpOGOYO �O}O�O�O�O�O�O$_ �O_Z_1_C_U_g_y_ �_a?�_�?�_�_2o	o oho?oQocouo�o�o �o�o�o�o) ;M�q���� �����_`��_)� ;������ޏ��Ǐُ &����\�3�E���i� {���ڟ��ß���� F��/�A���e�w�M� _�q���������� +�=�O���s���ҿ�� ��Ϳ߿��P�'�9� ��]�oρϓϥϷ�� ����:�կ��'ߔ� �}ߏߡ߳������ ��H��1�C�U�g�y� ������������	� �-�z�Q�c���K�]� ����
����R) ;�_q���� ��<%rI [m������ &/������/%/�i/ {/�/�/�/�/�/�/�/ ??/?|?S?e?�?�? �?�?�?�?�?0OOO fO=OOOaO7/�O[/�O �OqO�O�O>__'_t_ K_]_o_�_�_�_�_�_ �_(o�_o#o5oGoYo �o}o�o�o�o�o�o�O 6�O�o~Ug� ������2�	� �h�?�Q���u����� 揽�Ϗ���R�)��;�M�f��$DCS�S_PSTAT �������Q   t�佐ɐПԐ  �Ν (�  �x���͚���ԟ;�� W� t���k�損�����e�����¯p�������SETUP 	��B�x�k�� �4���U�D�y�h������T1SC 2
4�f�m�Czk�ݿ��ͺ�CP RȼD�D.L�^�  �ϔϦ�u������� ���$�6��Z�l�;� }ߢߴ߃���������  �2�D��h�z��[� ���������
���.� @�R�!�v�����i��� ��������<N `h�8ύ�&�� ��/�Se wF������ �/+/=//a/s/�/ T/�/�/�/�/�/?�/ �/9?K??o?�?�?b? �?�?�?�?�?O#O�? GOYO(O}O�O�Op�O �O�OpO__1_ _U_ g_y_H_�_�_~_�_�_ �_�_o-o?oocouo �oVo�o�o�o�o�o �o);Mq�� d������� �I�[�*������r� Ǐُ돺O�!�3��� W�i�{�J�������՟ ���ȟ�/�A��e� w���X����������� �֯+�=�O��s��� ��f���Ϳ߿���� �9�K�]�,ρϓϥ� t������ϼ��#�5� �Y�k���Lߡ߳߂� ���������1�C�� g�y��Z������� ��	���-�?�Q� �u� ����h��������� ��;M_.�� �v����% �I[m<ߑ�� <����!/3/E/ /i/{/J/\/�/�/�/ �/�/?�//?A?S?"? w?�?�?j?�?�?�?�? OO�?=OOOaO0O�O �O�OxO�O�O�O�O_ '_�OK_]_o_>_�_�_ �_��_�_�_�_#o5o Gooko}oLo�o�o�o �o�o�o�o1CU $y�Zl��� �	���?�Q�c�2� ������z�ϏᏰ�� �)���M�_�q�@��� ������ݟ���_%� 7����m��N����� ǯ������ޯ3�E� W�&�{���\���ÿտ �������A�S�e� 4ωϛ�j�|����ϲ� ��+���O�a�s�B� �ߩ߻ߊ���������'�9���$DCS�S_TCPMAP  ���g��Q @ U����w������	�
������� � ��������T�����U��� �U!�"�#�$�U%�&�'�(�U)�*�+�,�U-�.�/�0�U1�2�3�4�U5�6�7�8�U9�:�;�<�U=�>�?�@W�UIRO 2g��x������ �������� 2D Vhz�����������3E Wi{����� ��////A/S/e/ ��/�/�/�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?|/O �/9OKO]OoO�O�O�O �O�O�O�O�O_#_5_�G_Y_k_}_O�_S�U�IZN 2g�	 �x�v��_�_o ��_4oFoXoo|o�o �ooo�o�o�o�o 0�oTfx;�� �������>� P��t�������m�Ώ ������(�:���^� p���Q�����ʟ���  ���6�H�Z��/� ����q�Ưدꯩ_Z�UFRM Rf����8�@�R�� v���c���������� Ͽ�*��N�`�;τ� ��qϺ��ϧ����� +�8�J���n߀�[ߤ� �ߑ��������"��� F�X�3�i���{��� ������#�0�B��� f�x�S����������� ����,Pb= ��s���� �(:�^pK� ������/$/ �H/Z/5/~/�/k/�/ �/�/�/�/
?2?D? ?h?z?U?�?�?�?�? �?�?
OO�?@ORO-O vO�OcO�O�O�O�O�O ??*_<_�O`_r_M_ �_�_�_�_�_�_oo �_8oJo%ono�o[o�o �o�o�o�o�o_"4 �oXjE��{� ������B�T� /�x���e�������� ���,�ˏP�b�=� ����s���Ο����� ��:�L�'�p���]� ������ܯ�ȧ