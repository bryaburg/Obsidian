��   X�A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����CIPS_C�FG_T   �0 $INTE�RFACE  �$DUMMY1�B2B3B&SE�T/ @ $�MODA8 _S�IZ}OUT�DATE_FIX~�CSI_VRC �    ��$$CLASS ? �������O��O� VERS�ION�  �Z�$'1 �O� �m @r �
��� �0�  -@