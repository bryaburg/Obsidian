��   !��A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG� ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S�ETHOST� � NSS* 8��D�FACE_�NUM? $DBG_LEVEL��OM_NAM� �!�* D �$PRIMAR�_IG !$AL�TERN1�<W?AIT_TIA �� FT� =@� LOG_8	��CMO>$DN�LD_FI:�S�UBDIRCAPė����8 . �4� H�ADD�RTYP�H N�GTH����z +LS�&�$ROBOT2P�EER2� MAS�K4MRU~OM�GDEV��PI�NFO� $�$$XC�RC�MT A$x| ��QSIZ��X�� TATUS�WMAILSER�V $PLAN~� <$LIN�<$CLU���<�$TO�P$CC��&FR�&�JEC��!�%ENB ^� ALAR�!B��TP�/3�V8 S���$VAR79M� ON,6��,6APPL,6PA� -5B N+7POR��#_1>2ALERT�&�2URL }�3�ATTAC��0ERR_THRO�3�US�9�!�8R0CH�- YDMAXNS�_�1�1AMO	D�2AI� o 2A� �(1APWD  �� LA �0�ND�)ATRYsFDEL�A�C2@�'`AERS�I�1A�'RO�IC�LK�HMt0�'� X�ML+ \3SGFReM�3T� XOU�3fZ G_��COPc1V�3Q�'C�2-5R_AU�� � XRN1�oUPDXPCO�U�!SFO 2 
$V~Wo�@�YACC�H�QSN}AE$UMMY1�W�2R"�RDM*	>T $DIS���SMB�
 T M�	BCl@DCI�2AI&P6EXsPS�!�PAR�� `RANe@  ���QCL�� <(C�0�SPsTM
U� PWR��-hCfSMoC l5��!�"%�7�Y�P�% 0�fR��0�eP� _DLVH�De\aNo3 �
j�hX_!`�#Z_�INDE,C_pOFYF� ~URnyD��*s�   ts �!pMON�r�sD��rHOU�#�EyA�v�q�v�q�vL�OCA� Y$Nާ0H_HE��rPI"/  d	`GARP�&�1F�#W_~ �I!Fap;�FA�D�01#�HO�_� �R�2P$`�S�wTEL	% P dK  !�0WO�`� �QE� LV��k�2H#ICEدڀ���$d�  ��������
���
��`S$Q���  �Zc�$'0 �
����F����"�S�L���$� 24� T"�����e��� 4����! �ʟ����-�4�Ɵ��8�I�L����p_V`4�� S�z�������¯ԯ毀��
��.�@��� _?FLTR  �?�W �������!�ޛnx4�2ޛ8�{SHE`D 14�E P'��I�ٿ ��:���^�!ς�E� ��iϷ��ϟ� ���$� ��H��l�/�Aߢ�e� �߉��߭������D� �h�+��O��s�� ����
���.���R�� ^�9�����o������� ����<��r5 �Y�}��� �8�\�Cy�������PP�P_L�A1e�x/!1.9"0/��8%1I/�2551.�%@/��Q�7#2>/P.� d/v/�/�/�&3�/P.-0�/�/ ??�&4.?P.�0T?f?x?�?�&5�?P.@�?�?�?O�&6OP.�@�DOVOhOzOT�aP���t(�{��Ӱ��� OQ� ��N<0_ e_w_J_�_�_�_�_�_�_�P�_%o7oIoo moo�o�obo�o�o�o��N�o�T�5 |�
ZDT Status�oD�����}iRCon�nect: ir�c�t//alertb~���+��wt�Y�k�}��������2A�d�RJ������  ��$�6�H�Z�l�~��������ƟQs$$c�962b37a-�1ac0-eb2�a-f1c7-8�c6eb571d?066  (H��@l=�O�a�s���A
��X�'R��)z��`P��*s,P!T,$4� 񯨰*!߯��@�'� M�v�]�������п�� ��ۿ����N�5�r�4Y�����&%P7DM_Q	&+"?SMB 
&%U��#l��O���� �I�ff|������_CLNT �2&)9�4+t 	�|�#|j߯ߎߠ��� ��������Q�0�u�f������
.S�MTP_CTRL' R� P%��4� 	t��"�c���R���v�H��#|��N�Q�����7������ ��USTOM' ���&P� �TTCPIP����'xU"R�i EL$&%#Q�> H!TP	���rj3_tp�т��+ ��!K�CL�������!CRT.uR��!CONS�v�
�ib_s'mon~r