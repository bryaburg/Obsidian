��  	��A��*SYST�EM*��V9.1�0170 9/�18/2019 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ���AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP�fBI�IZ@P�_�ALRM_RwECO"  � wALM�"ENB����&ON�!� MD�G/ 0 $?DEBUG1A�"d�$3AO� ."��!_IF� |�� ENABL@�C#� P dC#U5K��!MA�B �"�
�� OG�f 0CU�RR_D1P $Q3L�IN@S1I4$�"PPINFOEQ/� �L A �?1~5/ H ��79EQUIP� 2�0NAM�� ��2_OVR��$VERSI�� � ~0COUP�LE,   $��!PPV1CES0��!H1�3�2> �1�	 � $SO{FT�T_IDB�TOTAL_EQ2� Q1Q@NOTBU �SPI_INDE�]iEXBSCRE�EN_�4BSI�G�0OKK@P�K_FI0	�$THKY�GPA�NE\D � DU/MMY1d�D�!R�E4�A�RG1R��
 � $TIT1d ��� +Td�+T� +TP+T5)V6�)V7)V8)V9)W0 )W2W�A+UFW
Q+UZW1dW1nW1xW 4V��R�1SBN_CF��!�0$!J� ; 
2�1_CMN�T�$FLAG�S]�CHE"=$Bb_OPT�2 �� ELLSETU�P  `�0HYO�0 PRZ1%oc�MACRO{bREPR�hD0D+h@�؞b{�eHM MN�B
1�0UTOB� U�0 }9DEVIC(STI�0�� D@13��`BEdf"VAL��#ISP_UNI�p_DOv7=yFR_F�@K%D13��/A�c�C_WAx3t�awzOFF_�0]N�DEL�xLF0pq�A�q�b?q��p�C?�`�A�E��C#�s�ATB�t���MO� �sE 	� [M�s��&�wREV�BIL:���XI� �R 7 � ODq`^��$NO`M@���0V�l�/�"@i�� w����1X�@}Dd p E �RD_EV��$�FSSB�&K`KBoD_SE&uAG� G�2 "_��B�� V�t:5`ˁEC�0��a_EDu � �� C2�}`S̄p�4%$l �t$�OP�@EB�qm�_�OKԂUS�1P_�C� m��d\�U �`LACI�!�a����<� :qCOMM� �0$D��Ñt@�pL���O�B6�IGALL;OW� (KD2:�2�@VAR)�d!�|AB 6�LO@S �C ,K>qA�<`Swp�N@M_O]n��w�CFd X�0�GR�0��M�N�FLI���/@UI�RE�84�"� SW�IT=$/0_Nc`S��"CF_�G�� �A0WARNM0lp�d�`LI�J`wNST� COR-��bFLTR�T�RAT T�`� $ACC�aG�� L�>r$ORI�.&vǧRT�`_SFg��`CHGV0I��d�T��DA�Iu�T·���� �� �#4aԂ�HSDR�B�2�BJ; ��C���3��4��5*��6��7��8��  f�z�l@�2� @� TRQB��$f��ʀ���c_U�����0COc <� ������x3�2��LLECA�}!�MULTIV4��"��A
2FS٠I�LD8��c� DET}_%b  4� STY2�b(�=4��)2(���08԰�� 
7$��"p��*�a=`�* P�TO��:�E��EXT����p���B�ђ22��,:��@��%b�.'�B �;�E� �"E�/%ua��L� �3s�9�I� Gғ؈/A�Ƌ�M�� �� 7ՋC�! L@�0U�� LׯpA²$JOB6�����Ǳv��IGC�" dǀ �����L�-'l��;��ƧY��`��b# t2ǀF� �CNG�AiBA� Ñ�����/1������0����R0��P�#p��6��$��@p��t6q:Q�
2JQ�S_RB�qCTJT�TYtJ3�D/5C�	@�ǧ��@� ��P��O'л!% \�0RaO�6� �IT}s� NOM_,pn#`�c��ՠTU�@MP� � ��&P��� ǨP�	ѭ��RAl@n �3�5����
$TF'%#D3� T��kpU�1'�q�e%aHr�T1�E����ң�#Ѥ�%8ӢQ`YNT�"� �DBGDE�!'8�Q�PU���@ȟֽ�"��AX��"�uT�AI&sBUFφ=9t1#�1( �װD&�J`PI84'aP��'M�(M�)6 �&F>�'SIMQS�@NwKEE3PAT��nЍ,"�"�MCb��)G�$��`JB��ĲaDEC[:� [5������* �I�CHNS_EMP��G$G��7�_�<�c/�1_FP�TC�6S���5�`��4�q y�V�x�K�x�JR����SEGFRAe�OUaP�T_LIN�?CP�VF�A���`�7$+ ���c_BNu�DBnr[�|�@*,` +� Ȧ9��A�0��AX0c`�5r�D���IX1SIZ\����D�FT�C�Z%Y�ARSa��CD@��IW\%@WX�00@Lp����0�VCRCӥ�sCCw��U%@�X�1խ�2�Mdq�U�1T��XxQ�UDѤ̣�YC k�p���4?`рf��FhEVFf�F\a_
�5F�0N�ftPX1��h��)�^Cq�+��VSCAO��AH�f����1'��-հy	��{MARG��D�U�F4@���1DWQ��r�0LEW�!�@�R�P0Ҹo�l�R��.� ���ϻ�����%ΡR� HANC��$LG)��a� ǐ��̀:��AY���u0RMr�3�s�����s4 �xRA���sA�Z�0E�B`�O��F#CT�gp�FԠ�R��0D0V ADI��O �����������)�)����SO�[���'BMPIDPY �1���AES7P^c��W
��N S!�B����_/  �PI,d?��40��b@_C�$�m�K�"U0ϑU:��1�TITq0�bV�%97A."Z_`.G2 ��� �!��vNO_HEADE��!~�w�l�0��z�S+�q�R9�����43 T��b�5C�IRTR�0�W�XLdMt dC�gRJ��{ ��!ERRLX�b �4�Q͠OR�B�$ᢳ�����UN�_O�p�P$SYASР4�͠��U��EV�J@�@DBP�XWOyP �5z��$SKc�"�aDB]T�pTRL��6̐��P�����IND&I DJ�d�_�`�!�������PL�A�S2WAzⰰE��D�!��!R\��UOMMY9��1Л |�DBO���7�E��!PR~Q 
pC���-���8 ж�$f�$Q�5�L�9+ώ���P �:Qώt��PC��;p�c�EN5E70Tq<��cþ��RECORj�=�H aO��78$L��9$Þ"�9���F@t�JA �_D�ʁ� ROS �"SK���rj�ׂ� 1���C�PA��>JBE�TURNA��SMR��U �CR�E�WM8B
0GNA9LJ �"$LA� ���:$P�P;3$Pj�g�<��!b�PC���PDOR@�Q����R�GO_3AW�"�MO���p� �ǠCSSp�STCY��>����0Ls�<�ID���2?�2M�N��OB�>&��j`I� ? P7 $@�RB�Bt��PIM�PO��I_#BY ����TJR&��HNDGj�@ �H�`�1���0{�DSBL=��s�N�0q�%�LS��A��0� f,�FB[��FE�@@��N�&�)0B? �$DO�1�C�pMC�0��I�4���R�H��W/ ?(ELAE�u
r;����Cq�s$^�q�INK�)[�UV�L��HA�]�QoP$|#oPp��(��� D �i��MDL 2C Α5��C���JoR�oR���	��g��	��[��'�SLAVrElBING ��#8��&�C�FP�@P` �p��q�������ouС�O!���!��ID�������W��N3TV�#�VE�$СSKI��`A�C/3	'	2IB�1J�f�1���4�SAFJ�C'_SV>*�EXCLUs����LrONL�0k#Y���s����HI_V�ɀ�RPPLY��Rb7sH� ~�#_M�b}# VRFY_��z�"Mas$IOj0����&��1IB�$##O����%LSR���4�Ǳ2N�.@a�P�-�$,��&AH CN�f@�a5N�F3t��GCHD�s�_�L�E &*�CP��4TǱ�8jŀX� G��H��TAn���!� w��hNOC
tIHlB�pTQоA ~7�D���$�I D� $��6�L-:C!qPCF_\ �NLHLC@��E�@Kb2�J��q�0x$(Bn� I eSG�`� K �ΐCUR~ЛѰ���A#�0����(��H(��FANNUN��j5�CN��@�������YQ��$Z�@V@�EFРI��L� @�`FR��	$TOT�Ч��03��ձ(5��\PM+�NIBK�M6�R��RA���TDAY�LOA�D��䴧R�5���EFF_AXIJJ�N��ڱ�O`T�À�_��QqO2@P�`�6`BcE�Kce� Nh Qw1a����A$p&aqP 09Q�an� �a�ӯv�DU�Яu�^�CA QjR���n �,�IDLE_PW�Gs�e�-�V��V_��`� ���DIAG�_�R� 1$V��SEs�T}�6q � <zǰR���Q�V��@SWsq��Cp�`�1e� �O1aOHGe�aP�P�IR��B >��b�ᑠ�:P�r 6��x�R��u���e� �Qh 6`,�:uRQDMW�uMSG�6�A�x�uarLIFE��BSQ@��"Ns�=r|�HQq�=rC8�SC��@@�N�YՐ�F3LA�3QOV Ј��퐰�SUPPO$n��"��_��E���_X*����Z�W� ��q�	��XZ_A�Y2o�CF�T(�)�;u!N�9uQ� �vn@�BICTlS{ `# CACHC���ؒ`�Et#��y�SoUFFI�� ��.�b�6��A�wMSWɕT 8(PKEYIMAGf�TM���SU��BQ�J|g�@�OCVIE}p��U hBGLx�P�?� 	�Q��0ʔV2@��ST !��YpŤհŤ��PŤ`ŠEMAI�� =��Q���1FAU�LK�W��<�u�AXb�U�h�3TB>P
nXC�R����X��&��0���LDEBU. �  AT���a?Y< $y����S�`�`IT��BU!Fꗤꗋ�N�!wp'SUB����C�#�8z��q�SAV𵲲�7p��Yчp�  VP ������~t�_��ֵ��PL�OT0���cP�� M�v��2s�AX��S]P� X��M#$�_�Gs�
G�DYN�_�q�PZ <@`D����+��rM�b*T80Fg�%�0{DI�2EDT_{�$��Q[E� GƱxQ&�C����A��ҷQ\� �� %�nT�C_R��IK�rb��B_�=RM�^��NB�DSPe�B�P� ��IM���ѥ5B�B*pUy�ހg�`�M��IP�Bӱq����T!H��y��`T�q��sHS�~�BSC����`V�P�J��R�{_D4CONVW!AG4R䍐�֥�Fsq�"d~������qSC8r�T�MER�$BџFBCMP�#A�E�T ]C�FU&��DU��/�o e��]2CD���g�� M���NOa1�Q^2B�;��U;��UP�1=�C@J��1p�8�z���P_H *J�L ��0����>P��# ���1���Q���Q��a���-���7��8��9P��s�����1��1��U1��1��1
1
U1
1,
2:
2�����2��2��2��2�
2
2
2,
3J:
3��3����3��U3��3
3
3
�3,
4:��EXT-q�Q`�������������'_�,�FDR^taT��VC0�n�v�D!J�v�REMrUpF��OVMu�zj%As)TROVs)�DT���*MX�,I�Ns)���*qIND�� ��
�(	�v���G@���s� ��|�bqDFf�� RIV�0����G�EARu�IOYuKc"��N��Q8aW�S��q����Z_MCM\g�v�G�F߀U@Η�b ,H�ȱ?� �A���0rq�?�1E9p�1@�H���9"c�P!�P���)pRI�в�E�TUP2_ d �P��TDDЪa���T�@�1GE�A��B;AC��e T����
(�)"�%nS�����IFI�q����@�oEPTr�2LUI�4�f ��`_�{�UR�q۱�����JਰT1sV`IW$$�BS�@�?x�@J%�CO�?�b�VRT�yPx�$SHOUaJP�A�SSZ�m����$BG_`MQnMQ��MQx��MQ��FORC1�^�BDATA�ag�KFU�11�S2:Ӹ�D���ah |� N;AV}���@R��_ S���$VgISI0�SC}ģSE�07P�eV`O�a$a�B�B�A�`^f$PO�PI�q�FMR26%i C"S��b D!6�^fH'O?a?s?�&(I�:uc"_:>FpGIT_�A�TpM6|-??=DGCLF�u�DGDY'xj���DCG5��?|�0!M3��jy��i T��FSJ���k P���r6�v�$EX_�q�x�q1���࿂j�p3�{5�v�Gf��6%l �� ��SWٵONA�k�QTl�h%�GR&@f�U��BK�U��O1�  ��PO�`K�7���
�:7�M6PLOO��y�SM�`E���1� p_E m ����� �TERMr��n��?AORI�r��o���0SM_#Є����p��5�P�q줆|�UP��r�3 -�!rm�@���)�n`G.�@pELeTX�ҁ�FIo���њ0��Ʉ%�o�$UFR)�$`>�X�����`OT��Ɓ�TA,�W`��NST�PAT!��OPTHJL��E��8'��X�ART�b�pYp����REL���SHFT��ȑ���_"PR���� �$��X�q�aE P��Ӵ�SHI'��dUz�� O�AYLO�� �a���@�0-Rȑ�QR��ERV���BC� �����`�@�n�@RC�1R�ASY1M��R��WJk���� E�3���B�U�B������Yp��P��Ӱ���r�OR�MF[c�p��Jds�R�7�p�ǐ���a0 HA�PTIV�t�2MA8�������A!��A��qHO6Pvtu aԮ��E6`[`OCQ��U��1$OP0!dFѩ�9S_!$P�P_ T�R���OYUL�ȓe�@Rƕ��o��[De$PW�R 0IM��ĢR_�J���P�ۓX�UDp�2�0�x� v@�$HhE!�AD+DR&H��Gʒ-є"���7�RbMaw H�S��	a`Z�`nZ���Z���SE�alc��HS�MN�Bx`B�F"��(�$�OL�� }�%����RO�Pa��AND�_C��=�¡�Ć�R'OUP��Բ_�0�RU�ձ1�xb0��:� `:�h!;���:���:��yPxbA`B2��AV#ED5��E���Jc�y $�P��_D��X�-R��PRM_��R4�HTTP_�=�HMaz (H�OcBJ`�[D$&�LE������N`{ G� ��@�_�!�T��N�S԰���HK;RL��HIT糫� NP��al�N�%R�F)S�l��Gm�SS� $J�QUERY_FL�A��"�_WEBS;OCb�HW&^��Ma|U�w�INCPU���QOc�P��& p�%~�%�t��IOLNKB} �8�RI@�$S�L\b$INPUT_��$��t�n>a TP SL��
Ma~[ q����~��1IO��F_�AS�rQ@$Lf@"�fAH�a��o�`�@a�j��HY'p+ �� UOP�u� `� I&�"� "s��P����i��"��D�IP_sMEa�A� X� cIP"����_N
��r���qI�s�)!���SP[B��~PBPB�G�ѭ��PM���A�3 l�p{�TA��)�A6P㰔n����`U%��PST&BU�`ID�p��6P|%z�{%��$!w"����5*�h$I$| N�(�`�%�IRCA_CN� _ � �@�� CY��EA
1a <g��'7�C��=�~#�x�DAY_� (NTVA�E� k7�敜w#k7SCA��k7CLq�!-Q��"`�A���/�$��%�5N_�T�C�B� �"Y1�@� ��P`�A�� {!���_8�Q 2� �O $!iA�A�� q$RF�R LAB���pA�`vGUNI�dC̀ITYb$!&բ�R��
P�s��C�UI�URL�P�$A��EN?�ۡ�Q�����T��T_UA2 ��J �Q��$$R"�J�@ Ra$P"�`A��.QJ��9R#FL�pA0x`
MS5s�
�UJRIe� �� F�pq�P��yR=D�3$J7��RJ8�Y7�p^2�R�W�7uF�P8�Y�QAP�HIBpQ�S�WD��pJ7J8ڢ`L�_KE�@  ��KG LM�! 7� <�0XR�  �3WATCH_V�A�Ѱ��A�FIE�L��y��(b�u�� �`��V��V��aC�T�@�f����LD�M� x4��_�M��ΡD�1Q�LNsTK����COO���fNF��fTa�`�����JvP�(�����LG�d�� !~�)LG_SIZH�9�[uMRYw� ZvFDexIYxpxl�gv|x ��ZvWpf�`s�vop�v � �v�p�v���v�n�:P�_��_CM��#�Lg+�'�F$�1�K��Wp��(Vqc� bqp�opp�� p��p|�Io����pp��pp�Wp�RSK`א  (��0LN�Q���U��DE6�E�`�A����԰L���DAU"�EA��G 6��8�.�GH7������ BOOO���� C
�IT0��l�/RE* ��GSCRX��D��|��"�MARGI� �з���U�ᒍ��	S.��W������JGM�MNCHL�C�FNb�K@���@>�UFL���L�F�WDL�HL��STPL�VL��@L�s�L��RS��H��h��C�����A������U ��`�򗈃��`S�G0�	�POW�����`��,�6�!N�EX�TUI>�I�pC0��q.�ֳ�ֳ<��A@��o���������N�����ANA�+tAV�AI�P�Ա3�eDCAS\0b�R�p�R�OX�EOd�SA3��o�S{�֘IGNpp�0�s=���`*A[�DEV��LAL�aN �w"Cp��`�!Tr�$fw�H� 4dQ��A� �B���0b  ���+S1J�2J�3J�$a8��S�Cp� �@�p)t}��~|%�����r����Q��ST[R�9�Yr�� �$E��C�ۘP����p	�qa��Bq� L  �p.���e������j�a����_ � �������3��ޘ��MC���{ �� CLDP[>�eTRQLI�AV���FL!��lQ��b�1Dwa����LD������ORGQ��~�RESERV(�M�4M�?��lS� ��`�������#SV����TR	1��}��RCLMC���M�_���J ���OMDBG�Q�5`1sMA�dU0FC�%U�T8�r%E�P���MFRQL�� � KyH_RS_RU�b��DA0$�FREQ�6�u�$�YwOV�ERj �s���~VPnU�EFI� %G��D3u Yz�� \8P��T$U��Bg?�`�1PSI�9P	��`��D"���U� %?( 	ޜ!MISCkU� Yd����RQ7R	 �pU07P�鱎A�X�b#`��EXC#ES�BdQdM)@oQ���`u�di�dS}C�� � HA�_I@.0+��/ �MK�D��d�%B_�`FLIC�B�B��QUIRE� �pu+O�+�� L:d�M�E� ��{��� �b�c����ND�g0pP����Lx 3�D;�
�INAUT@��
�&p�P8��Nr��q��"s��!PST�LoQ� 4�0LO�C��RI�@��EX��6ANG*r.O[DA]�qrBzPbMF�b�u����c⽰m��5�$SU�Pv�W FX1PIG}G� � ��` c��q��c�
�c�@� ��5I��EH��TF5 t��0�TIl`C�L�1�IN� tV�0MD�AIB�)�FX��D���GH�0�Q�DGDIA�Q�C4PW�P�D0ѧ��ED@�)aqOjS��pP� �CUppV	P��.��Oؑ_ � �`{Еӿ3 4r��pB|XP|^r����PP{X�KE�T`e�-$B8� oV��ND2��Pc��Q2_TXl�XT�RAX��R���� L�O:���d"	 f�CR.f&cW��MRR2h��� -a�A�� ?d$CALI��u�GF�jg2F�RIN�b�nc<$Rx`SWq0���c��ABC�8�D_J�P{!.�A_�J3�f
�b1SPH� P.P�d�m3�m(HQ9�.#uJ��3u4n��O��IM��MCSKP��bt7�?�btJA�MQb|�uyu8�u�w�0_AZ��/q��qEL��.r��OC�MP�3���RTE�s e1�0pe��1���� �Z�ScMGՠ�@��JG���SCL��5SPH�_��M��f���.�u`RTER�`nc��k`_E���b A0ؐ��M��DI�qQ��23UdrDF`vāLWʈVEL���INx���_BL X�.��Yq/J�������IN���]`��CR9�ْ�28�6�_T �F�a���W �^�"�k���L�D�H��P\a���$aVw`3_���$=�X�~&�$��� �R6S]`�H ��$BEL�pm��_oACCE�� 	�<���IRC_��q�@�NT��$SPS���L`�0 M���9�.��1G�/��Q���$���3S�T@�_G�ؒ�����8�7_MG}DDء��~FW��@���$����DE�PPA�BN[�ROg�EE ˢK�B����qK� ��`$USE_tv`�P� CTR��Y4�ꐪ� ��YN�gA鰢�Rp�A��M:NQ=�ҠO�v�ϴINC(T�1������Yq�ENC��L��A.K���H�IN¿�IS�8ť@O�NT|��NT23_Ȃ~f�LOـ~|�� I� #��΀#$ ���h��#"CQ�M�MOSIݡ<"[P���MPERCH  ����� �Ǚ1��lA�� ��lA�w�r������Ps	AS�E�L��Ps7'Ow�N�@�ʄ֟�TRK��R�AY"c?�!�� S��ոӔ0�v!��P MOM鲎"C�HP$�jg�ӆ�g�T`�DUXp��S_BC?KLSH_CS�F� : �ƴ ��-e��o�|���uCLALMJ�p@�Њ���CHKep|�@�TGLRTYp@ �S8ėE5�A_�3��'_UM3��C3桸Z�� LMT�`_ALG��s%��A0�E*� K�=�)�@�F�@�p9�NҌ�)�PC��)�Hp@� ܥ��CMC�U\��CN_�bN�SL��;sSF���V����A.ǃ���S�/��CAT��SH�3�b�  ���/�/�eT�i�f٠PA���_P����_fpZ�����eq�����JG�0��Ӏ�OG����TORQU~��e���� �e"���� �B_W���@ّaʓ`Г`IhIvIГF�0S:rX�Iq�VC�0!%�1�ڠ��q��JRK�!"&<PD�BX�MtS<PM0_sDLʑ_�GRVg``$ʓ`$ГA!H_%c8?#���*COS�+�p�(LN# �+��$ʐ �)=��)��*�,�<%1Z� ��A!MY�!:8�"�Q�+[9THET=0��NK23Г�2lē� CB�6CBēCz`AS�A�2��1ʓ�1�6SBʓ�2�5'GTSkqZ�C�a����&�J�#$DU��h�6Bjb��EG�eQ%�_��xNEht�@I� �������y1�A}5�E�G�%�(�!LCPH�%�B^ńBS� �C�%�C�%�B6!SZ(6�@V�HV�H���LUV�JV�KV
[V[UV&[V4[VBYH�H@�F�R�Md�X�KH
[UH[H&[H4[HBY�O�LO�HOsi�NO��JO�KO
[O[O*&[O4[O(6F�B�1�y�%t�GSPBA?LANCE_J16s�LE�0H_}5SP�>��&^r�&^r�&PFULCbx�rqw�r�%�K�1��UTO_<����T1T2�y
�2N���V��tM��Ѡ�pi@Z��	�Tu�O����QINSEG���REV���G�gDIF��p�1�U�6��1���OBK���j#�2,V���I$L�CHWAR4���A�B��$MEC�H�1J0��ǁ��AX���Po����G���p�� 
�?�0�RO�B��CRM�#���)�  �C�_�T� � x $�WEIGH��w �$�C\�� I����I9Fv��LAG����qS��:���BIL��cOD�Ы�s�ST�"s�P:���t���N C�L��P�
������  2���x�D�EBU��L|�Ē�5@MMY9C�9�N8�$�w $D|� ��$�� l1 �$L�DO_:�AK�� <_�ޖ�p��$���@B����NJÁ��_���� ˒O�� ��� %�T�7�?��TL��F�TgICK����T1N�%֣=�ߠN���pu���R\ఱ��񥩂���U�PROMP��E~�B $IR"ற��8�X�w�MAIF ���Q�_��P�P��X���°RU COD��FU����ID_�����8�2�>pG_SwUFF� ��4��X��DO��/�������GR����Ѵ �ݴ��赩���-Ѵ�U�퐱_�H�_F�I�9G�ORDf�� R��36s��H®�N�$ZDT暵�ʒX��4{ *W�L_NA���ߠ���DEF_I �ȡ��������𦿔`��������ISm@@# m�|@�0�����D6�4���D�p(?�f��DO@pl�LOCKE�˳�`��2�Ѳ˰UMе ��Ѵ��Ѵ��Ѵ>�ݲ ��ܵ��ݴ�ݲ��2� 2�賴��赡���� �9�w�͸��P}� ���,т@F�W�ر�Ӟ6���TE��Y��� ��LOM�B_����0s�VI]S� ITYs�A�}O��A_FRI�s��~�SI,��naR�ܠ7��7�3��s�WB�W�Q �% _���EAS{����P| x�W�8�45�55��6|�ORMULA�_I��G�ǵ� h 
�7�C?OEFF_Oá&�H)á�0Go{�S���5�CA�p:�L�ˑG�Rm@ � � �$���rv�X��TM�ד��ɢ�ӭ��ERI�T�Ԑ�퐳�  �rLL�p�SΛA_SVk��$���퐴.0��퐵 ��SETU,�MEAG����t�ˑH�>L�� � (� ���lقl��Dw��ߠ�ќ�}Ԃ]d�����y��G�xг[@��P�R�EC[�qɑSKy_Apy� P_�?1_USER�q�2�$��*4 �qVEL@� ��-"!%��Iz��B��MT��CFG>��  �]�=OςNOREJ���~l"�OPWOR�@� �,B�SY�SBU�P�SOP(�!��T�*U�+X�1P��K"�%PA qX�#˂�OP�U����!}����� IM�AGz�� d�IM� 5IN���"3?RGOVRDfP�#	 �!P� 3 �|@g�hl�i5ЂL��BT:B>lPMC_E���!��N�`M�2��1����H1SL|p��{ �R�OVSL�S��DEX\���5a@��8_H0�7�I0��3��3GH�4CC�����5CAGI0_Z�ERl!�2:��O @ _C�O��RI����
�Fg��I��A�A��Z�EGA��� H_�̀ÐATU�Sk,�C_T31DX�FB� �F�ApV�p��C���� Dc� � �2�B�P-��AM�- �r1XE�@x9RMR�TvC�}@`��@UP�H�&�PX;�V�1��3�7R �PG�Y%�� $SUB��A�E��A�CJMP�WAIT�PC�UL+OWςFʡM��ЁRCVF_��ς�QKRE`F0���CF@�RLς�<gIGN�R_PL�CDBTeBÐP*�ЁBW�d2dt U��1eIG�!x!��qҀTNLN0f��bRT{3NO�N<!��3PEED�P�3HADOWÐ΃t ERVE�3�d�2�Q���SP�p � �L_�瀼��`1�tU!Nq��[p�QRTPNC�LYw���AP!P�H_PKTZ#�~b"RETRIE�C�x"�"+�VqD�FI�_r� �R�Zp�t �2�d DBGL�V@cLOGSIZ�܁�ZpaUm��tD\�c�`_TXτM��YC�B�EM�}R�s|��ˆCHECK~`p��`L �� 0@�vx9�ALE�Qx�P�A�Ў���SrIP4�b��
AR�r��N�=���@O��b��AT��xc��v�pل��1sUX� ZB��sPL��Z$� $d!~��SWITCH�r&E�WO��A����LLB��� /$BA�DvӞBAM�@.�C=��A�,�J5�`N!Y�6|_��_KNOWO�4u�L0U�AD/�c �
pD ��PAYL#OAq9ී_�A��T�!��Z��L�Aj���LCL_�  !4��S�?!�]2�F�C� ��p�� I��R� ��W�d@P�B��� _J@r�~�_J�� !SPTANDq��������Q��PL�AL_� ��
pA�BT�1��C�D��E���J3��Ŧ� T PDCK�0)Ҟ3COMH�PHգ��BE.��կ���X|a�0 � �\�`��D_1��2�DMAR@Q������|��:PRTIA4ùu5ù6�MOM��@ϳ�ܳ��V B`�ADϳ�ܳ��PUB�0R��@�ܳ@��:����� L$PI�4�at�!P��=Aܙ��I��I��I�à���\��ơQ���Q$RO�c���E�cHIG��ce �d4��de9`.`4�j��C�9aR�9aeSAMPHP=���4ק�eN��� &��� �� !"�ԡP���`���ٔ�!"R��ȴ�Տ�m���IN5����<�X�3��b>�~�U�~��GA�MM*�S�A���qGET!�FIO��c��>"
WIBF�bI<l�d�$HI���A�@!"�E;� �A�=�.�LW�[�R��=��.�X֚`ǡC�heCHKV0�@�F
�I_�Й�>"1� r�v�$������1����ţ �$�� �1���IRCH_D#��P$d�LE;!!�At^�< }ʧ`MSWFL3d�M��SCR�X75 2�p��O����F��ϰ���	�`��Pn�S�V#��P�pCUaR�#f�pSAA�Xn4A�NOb�C�A �c�A��r�ȟڟ�Ȁ�����������DO�aA���q���
� .ؚ">�^�j�?';%�����Mq�� � ���YL��r�$�����p�%�r�'@`�@	 �"�#r�(0� @a7Q'M_Wp�"�"`��#��s!MG`�+��'ġd�4���5�Rl�9M2wB� ��q� Έ4$WQ0�5ANGLa�Q0:�O2A�@O2H�O2�X`;�No�P�����sw�XGpOI��v�Z�5l�`r�� -���OM�� ����ư�pg^��rLb�_�R� | �HN﹛Fܳ�F:� NȺ�G�F����߀([�}D�߀�D�P���PMON_�QU�� � 8�:�QCOU:�Q�TH|`HO�"FPH�YS��EST�FPU�E1P7UpO�T� � gpP`�bRU�N_TO�#�PO!�� P���U!e�#INDE�sc�G�RA� ܀� 2� N�E_NO�T�UITxj �QsPINFO��er�[a�"��O�Ib� (��SLEQ%�.a�.`�V*ayS��p�� 4:��ENAB}2�PPTION���d�g�d�bcGCF�q� @b:�J0v�R����R�hhq�o�d�2��EwDIT� ��pR�0KE�&�$�E,�sNUwxAUT]uCOPYE�!�6|�iM�N@pD{���PRUTq2 GrNv�`OU �$G�R|�tyBRGADJq-�y�X_� I\�0(�v�0�vW�xP�x� ��v=ӻpBbN��_CcYC}2�p�qNSge9� w�LGO��(��NYQ_FREQ�W�W���\����SL�򐞂T��q곉�&�CcRE��QS��IF����SNA��%��_}GjSTATU�@<j�WMAIL�Ҁ�yIuATLAST偼�.�ELEMka�� ���vgFEASIxa?"��� � �&� JE��b!���I�P���S��IQPyz�AB$�a�E�PA�V���~�����X�U_�!�V���ǖRMS_TRt�v�g ��3^�Bb �Ɣ rP0��3�݊@	Q� 2� d�4R�7��� 6��.0 �!��b���NnDOU�SbN�c�0�PRd l`�5bG�RID�Q�cBAR�S%�TYycj� �O\
�q� �Q_���!�pݢ��O�0hd�� � � �@PO�R�S����SRV���)&��DI_T���?�R��\��\�4�Z�� \�6Z�7Z�8�>�zAF��ka�~P$VALU��47��QPF4��� !!teX�Q���1F�`AN3�́Rp|a�5�TOTAL��,�1A�PWI�I��W�REGENU�j��C�XӘ�Sa�Q�,PT1R��W�U�_S7��j��cV�q�d�¢b��E샩�KQ4��R,p�7V_HƠDA,C����S_Ye�2m�S�� AR,@2� >�rIG_SE����d���_�P��C_Ѧ�$CMPp7��DERtKБ�I��Z���\�Ba�0Fq0HAN=C2Q� p$�veq̂ ��INT=��g�0F�S�1MAS�KȃĐOVRQSP #P��H@��vầ�V������pb��V���Ѧ�OPSLGT�ka�`�=n��02?�H�S8�"����U��V�rP��TE�0İ����o��Jb�]}�IL_M|��w���@TQ,P��Q͐�j�"V2�C@�P_�VJ�Ma�V1`�VU1n�2}�2n�3}�3n�4}�4n�#���!"#�`���!"IN	VIB<0:�' !�.2*263*3
64*46p:���Np�T $�MC_FOPdB$ LBN��5�Mn1I�Ӳ~� �@5B���� KEEP_H/NADD�!����	C�1��ݡ���O%Q�zp�2 ���REM%@G� �JafU���eHPWD  ;�SBM���?COLLAB.4�h��3���`IT3���0UrNO5AFCAqLt2��4� ,7`�FLz0��$SY�N� ,M�@Co��~V�UP_DLYq=�~RDELA= H�ZɂYPAD,A��QSKIPS5� i���PO�0NT�!g P_�P�R�'�P �2g��'���)�a�)s� �*���*���*���*���*���*9�q�RA�hd� XJ�'���M}B3NFLIC�S�[0T�US����WNO�_H[ DHq�2IT��r<0_PA�PGN�� ����UҐ�W�`�6M���NGRLT= �Q�q�����8���1�T_J�!�6�BbAP��WEIG=H�SJ4CHxP�4cOR��4$�OO+����d��6J	���A0aA��nCIHOB`�`��:�J2s0q�pcX��TV��A�Q5��A�p`��A�Q��1DC���� �
pR�cR0P9�R���JIR�B9�RGE�`c��C��FLG�p�PH�d9��SPC�S�UM_|�@��2TH2N���_@�A 1� ��s0ݡ4� �� D����I��2_Pd2�SS����]�_L10_C{�� ܑU�� ��p$ �P2�Y��C�;�� a�D��aZ��Q�C�7c���hқ�NK��V�МP� P��D�ESIG�RV�VL�1�Y1�VTcg10a_DS��	���vOp11q� l� `��!��ATCp�t��_��bIND�����aOp9��b�2HwOMEr ��d2�b��o�o�o	(-a �d3�b�Pb0t��� ;0�b4�b�������'�  �$$Czh�SBP���ā�77 ��	�S�I"�π��Z�$AAVM_WRK 2 ą� ?0  �5ˁ�r%��H� H�A	k�\��7ŀ�m�������[�Νڟj�`���'�/��BS�`��A 1�� <�t����� ����ί����(� :�L�^�p��������� ʿܿ� ��$�6�H� Z�l�~ϐϢϴ����� ����� �2�D�V�h� zߌߞ߰��������� 
��.�@�R�d�v���?�C( AXLMT�BP���X�  dƝ�IN����PREoPE������_�C_��O  ��� c��� �ID �?ą��  8�d�^�p��������� ������9�-a���LJ��UPb��4�  �IOCN�V_lP�� ȴ�P�}�0��T�>�V@�  �1 �P $��`�����ŀ?�L �@ $6HZl ~������� / /2/D/V/h/z/�/ �/�/�/�/�/�/
?? .?@?R?d?v?�?�?�? �?�?�?�?OO*O<O NO`OrO�O�O�O�O�O �O�O__&_8_J_\_ n_�_�_�_�_�_�_�_ �_o"o4oFoXojo|o �o�o�o�o�o�o�o 0BTfx�� �������,� >�P�b�t��������� Ώ�����(�:�L� ^�p���������ʟܟ � ��$�6�H�Z�l� ~�������Ưد��� � �2�D�V�h�z��������¿Կ潝�LA�RMRECOV �M�����LM_DG -� �L>�_IF ����dFIL�E-066 UD�1 Ins Ge�neral��is�k 234 1 �mode J1 �at EOAT �chg,G1,A�1) 11��  uted VPL ���������!�3�W�w, 
< BA����8 �ߍ�AUT�O�� WORLD�o������ R&UP�PROGRAM �LLET_RIG�H����ABORT�E��QNGTOL�  �	 A� �Z�h��PPI�NFO H�� Gƞ������}�  T����-���-� �Q�;�M���q������������+� 1CUgy�������3�PPLI�CATION ?}������HandlingTool��� 
V9.10�P/23z��
16677557~H745891�цG264H=O�7DF1C���N�one�FR=A� 0��_ACTIVE�s  R�  #.��MOD ]�P��%CHGAPON�L?/c�V OUPLv�1p�� � �/�/�/
+CUREoQ 1	p�  ��,�,	?$5 94.��/??+?=?O?�a?�?�?.�N�"�%�4���"�:HTTHKY�?�?�?�?�?4OFO XOjO|O�O�O�O_�O �O�O__0_B_T_f_ x_�_�_�_o�_�_�_ oo,o>oPoboto�o �o�o�o�o�o (:L^p���  ������$�6� H�Z�l�~�������Ə ؏��� �2�D�V� h�z�������ԟ� �
��.�@�R�d�v� ��������Я� �� �*�<�N�`�r����� 𿺿̿޿����&� 8�J�\�nπϒ��϶������������%TO�C�/1#DO_CL�EAN`/$��NMw  H� �/�����	��-��.DS�PDRYR��%H	I= ��@�ߙ��� ��������)�;�M�8_�q�(MAX~�7��o'��X~Ԏ�"|�"PLUGG~ �׋#/%PRCP�B�������z���Ox��Y�k�SEGFW K5GR���ߙ����LLAP v��35GYk} �������/>R#TOTAL�����R#USENUv + d�h/�� RGDISPMMCU e��C]��@@k⒃$Ot���a#_�STRING 1�
O+
�M�H S*
�!_I�TEM1�&  n -
??.?@?R?d?v? �?�?�?�?�?�?�?O�O*O<ONO`OI�/O SIGNA�L�%Tryout Mode�%�Inp�@Sim�ulated�!�Out�LOV�ERRs� = 1�00�"In c�ycl�E�!Prog Abor�C��!�DStatu�s�#	Heart�beat�'MH� Faul0W9SAlerCYsOa_s_�_��_�_�_�_�_�_o z��+z��/oTo foxo�o�o�o�o�o�o �o,>Pbt8��oWORU �+ �qDo��
��.�@� R�d�v���������Џ�����*�<�N�PO�+$Qt��{]��� ����͟ߟ���'� 9�K�]�o���������pɯۯ�o�DEVw� ����?�Q�c�u��� ������Ͽ���π)�;�M�_�qσϕ�PALT0m����� ������,�>�P�b� t߆ߘߪ߼�������p��(��GRI�� �+`���:����� ��������*�<�N� `�r�����������N�F R0mx���,> Pbt����� ��(:L^<p��PREG�Ω ����//*/ </N/`/r/�/�/�/�/��/�/�/??vM�$�ARG_�pD ?�	���W1��  	�$vF	[k8]�k7�vG�9J0SBN_CONFIG�@�W;�A�B�1�1C�II_SAVE � vD�1�3J0TC�ELLSETUP� W:%  O�ME_IOvMvL%?MOV_H@$O�*OREPuO@:U�TOBACK�1�W9�2FRA:\� �O��0�'`P��H�� �K�0 �18/07/10o 22:%P18��8�6_H_u_l_�L���_�_�_�_�_oo���_DoVohozo �o�o)o�o�o�o�o
 .�oRdv�� �7�����*�\<� �  �A_�C�_\ATBCKC�TL.TMP DATE.D�̃���p����ˏ�CINI����E�6�CMESSAG�0��1_0�3�1>��ODE_D@�6��$�O�,��CPwAUS�� !�W;� , 	���0�� ��k���
����!����x|���=(�,		��W5 ��Ɨ���П���� @�*�d�N�`��������̩_�i�TSK  �o��A�1��JUP3DT#��d9�Z��XWZD_ENB8脸:B�STA�W1�9�I1XIS�0UNOT 2W5�1�0�� 	 ={�����pP�����}���eӖ�� �
Z	 x� �L�  #� .5 3q�����	�̱�h� �<�+= �"U&R�	Ϳ���
�4����\}π�MET 2���3 P��H��HY�|H9�{E�#UHS��AH�%;��@��|C?Nl�?��<�TN>����?���S�CRDCFG 1�W5�A ��5�2m�A�S�e�w��ߛ��O�U�9.��� ���!�3�E��i��� ����������N��B7�AGR��-�M�&��^�NA>@V;	ܘD#�_ED�1z��I��%-d�EDT-�RJ���� ��E��B�����2�_����D ����29����<����b�&�J��3QK�` R���.������4�A/ew�@e/�,I��/V	5�/ /�/1/w�/1?x/�/ ?�/��6i?�/�?�/ w�?�?D?V?�?z?��75O�?�O�?w^O�O O"O�OFO��8_uN_���*_�_�O�O�__��9�_=_oa_��_ao�_�_Po�_��CR8pO�o�o�M �o+ro�o�o&�s�?NO_DEL2�$��GE_UNUSE�0�"�IGALLO�W 1V�  � (*SYS�TEM*�	$SERV_GRj���pi�REG�uq$���pNUM�<8�&�PMU�pşLAY���PMPAL6�CYC10r~ⅎo�s���ULS���l����i��sL�����BOXORI��CUR_�&��PMCNVa���10��M�T4D�LIM����	*P�ROGRA�tPG_MIs������AL}�������B�ڟ�~$FLUI_RESU����
��C|C`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠ�x&��LAL_OUT ��{E�WD_�ABOR����I�TR_RTN  ���=�
�NONgSTOj�5� �x�CE_RIA_IL�p5�~�A�h�FCFG V�t~�u���_PA���GP 1����������ۯC�  >�@ࠪ@�@�@�@�Ȫ@��@��@��@���@��  D��D�|�|�8�S��@�@��@��@���|���D� D�|� ���pD3��=r|�F��j�DY���?��h�HE`pON�FIU����G_Pv-�1�� }u V�8�J�\�n�������|����KPAUS��1�~� �� ��	����|����s�����ݍ��b�� x��Ϻ�0� Z@j�v�� ���� DV�h�M*�NFO 1���� �� 	�ߝ�Ћ������XS����ؾ���@h�ፏ1k� D�z�?��EC2�������FB_�h��h�O�������!LLECT_���y� �9'E�N}�5��U"!ND-EA#I'�s>r�1234567890�'9b�q�ҧ/��&.c
 H��.c) �/?�l�/?^?;? M?�?q?�?�?�?�?�? �?6OOO%O~OIO[O mO�O�O�O�O_�O�O �OV_!_3_E_�_�ͅ$6�q2I+ ��X+>�"IO  �)U!.g4�o.o@oRo�W[TR��2!�](��bi
{_`n��"�]x�j��]&_MOR�R�#�� ?� 9B����u�y+�O=s�{�b���Q$
�m,��?����W��qR��K�ty���P"	&I/�����.�@��t�
�r�/'���ei@���|��cu ��a�hPDB�p�(�̉Tcpmi�dbg���1�*�:	�^��p�]�(�����^���l�`o���K��m��ƟCmgڟ3�����f"��{�<���Pud1�:��ɯ�j�DEFg '4c)���cّbuf.tx�tԯ"�կ��_MC�c)���Sdg�H��d�*V���ԕ���3�ˊC� B�!�C�9CaC��A֨lC2��IC�2�D��n�D��MD�9�CL~	D�mES�4��F,��F� �F�iE����
�Gb�7�kr S uD��w,�\rЪ��cĽ���`�Z�c�`x��,۱��Cf@�z�����^�D��E�H��D��D{�F���3ES�F�I3���F��E��}E{�H�F{��G�����  �>�3��C�r��n8�ѧ���5��ᧁ�cr��A�q7�=L��<#��ea��X����@�RSMOFS�T %�X��P�_T1w�DE -����a;���;�Q�s�m�?����<�M<�T�EST�+��R�C"./vC��A%�7�����?ї�aB�લ����C�������:d�T�b[�I�#/e�?��ʡr0�m�$r�RT�_�PROG ���m�%3�S�X��PNUSER  r%���f�KEY_TB�L  ����	
��� !"�#$%&'()*�+,-./�':;�<=>?@ABC��GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����-���͓��������������������������������������������������?�������Q'��LCKq�m�h�q�S�TAT�Y�_AU_TO_DOo&l��INDj$�8!QR����"-24:�!# STO� � TRL)�LET�Eo'{_SCR�EEN �j_kcsc"Ul�MMENU 11� <B�A�	/ X��/G/��$/J/�/ Z/l/�/�/�/�/�/�/ �/7?? ?m?D?V?�? z?�?�?�?�?�?!O�? 
OWO.O@OfO�OvO�O �O�O�O_�O�O_S_ *_<_�_`_r_�_�_�_ �_o�_�_=oo&oso Jo\o�o�o�o�o�o�o �o'�o6oFX �|�����#� ��Y�0�B���f�x����׏��������_?MANUALp�ZCD��2�ل���R��gߗ�?|(��g�L�@�3F� �B��7�z��7�0���$DBCORI�G��	�_ERRML/�4V�����>�P�b� �NU'MLI*�Wg�m��
�PXWORK 15V�-�¯ԯ����
�[�DBTB_� 6���b��t���DB_A�WAY��GC�P m�= �^�_A!L*��^��Yo�pm�&`�� 17��_ , 
���Se�(�v���a��ݾ�#�_M�I��l�@@�4�ON�TIM��m�ɼTƪ�
����MO�TNENDu���R�ECORD 1=�9� �"�#�G��O�����#�m�XE?CUTINGR�&� 8�J���T�{��ϟ�� ��������]���� ��H�l�~���ߴ�� 5���Y�� �2���V� A�����������k� ��
y�.��Rdv #��?� *�N�r�� ���;�_/� 8/J/\/n/��//�/ %/�/�/�/?/4?�/ -?�/|?�?�?�?!?�? E?�?i?O0OBOTO�? xOcO�?�OO�O�O�O�eO)�TOLERE�NCk�Bȴ�y�L����CSS_C�NSTCY 2>J���a�_���l_ z_�_�_�_�_�_�_�_ 
oo.oDoRodovo�o�o�o�oGTDEVI�CE 2?W[ F�#5GYk�}����#�HSHNDGD @W[Ƨ�Cz�z��JQLS 2A�m�G�Y��k�}��������IRPARAM BY��k�v�5��RBT �2D��8�<<ذ C;P���ª  �;P�Q��@W�F�E�?�d
�Q�HZ�Ԑ�\^���@��F�xM�+C�J��8P V�͐0ŌU��;�B�J�6U�ŅD�@����;�@��h��\�X�ńc�� ņ���Z�l�~����� ���د�7�� �2��ŅC�,�D
�D�0N�� 	��9�M<A�+�A���,A���A�?�A�U2Ŋ��YCs���B���4δ��Ō���|%Bw�q�B�0NB���QB�>_C�񹴿ƿؿ����? ��� gp� ~�H�ō-�O�a� ��I�wωϛϭϿ�� ����B��+�=�O�a� s��ߗߩ��������� ��'�t�K�]��� 7�������
���.�� R�=�v���cϑ���� ��������<% 7�[m���� ���8!nE W�{���g�/ �4/F/1/j/U/�/y/ �/������/��/�/ B??+?x?O?a?s?�? �?�?�?�?�?,OOO 'O9OKO]O�O�O�O�O �O�O�O(_�/L_7_p_ [_�_�_�_�_�_�_�/ �O	_6o�Oo1oCoUo go�o�o�o�o�o�o�o �o	h?Q�u �������� R�d��_��s�����Џ �����*�o3�E� r�I�[��������� ǟٟ&����\�3�E� W���{���گ��ï� ����X�/�A���	� ��Ŀ���ӿ���0� �T�f�A�o����υ� ���ϻ��������� b�9�Kߘ�o߁ߓߥ� ���������L�#�5� G�Y�k�}���E����� ��$��H�3�l�W��� ��}ϫ�������  ��	V-?Qcu ����
�� );�_q�� ��/��*//N/9/�K/�/o/�/�/�/���$DCSS_SL�AVE E�����!�~�*_4D  �.~3CFG F�%�3�dM�C:\� L%04d.CSV�/�{?�  ��A �3CH�0z��/g>�?��?�  �g6���1O�9A� J#(C�;g4��0��7,4RC_OUT� G�+OB�/_�C_FSI ?~�) :K g6�O�O�O�O�O__ F_A_S_e_�_�_�_�_ �_�_�_�_oo+o=o foaoso�o�o�o�o�o �o�o>9K] �������� ��#�5�^�Y�k�}� ������ŏ����� 6�1�C�U�~�y����� Ɵ��ӟ��	��-� V�Q�c�u��������� ����.�)�;�M� v�q���������˿ݿ ���%�N�I�[�m� �ϑϣϵ��������� &�!�3�E�n�i�{ߍ� �߱����������� F�A�S�e����� ����������+�=� f�a�s����������� ����>9K] �������� #5^Yk} �������/ 6/1/C/U/~/y/�/�/ �/�/�/�/?	??-? V?Q?c?u?�?�?�?�? �?�?�?O.O)O;OMO vOqO�O�O�O�O�O�O ___%_N_I_[_m_ �_�_�_�_�_�_�_�_ &o!o3oEonoio{o�o �o�o�o�o�o�o FASe���� ������+�=� f�a�s���������͏ �����>�9�K�]� ��������Οɟ۟� ��#�5�^�Y�k�}� ������ů����� 6�1�C�U�~�y����� ƿ��ӿ��	��-� V�Q�c�uϞϙϫϽ� �������.�)�;�M� v�q߃ߕ߾߹����������$DCS�_C_FSO ?����?� P � �\��������� ������"�4�]�X� j�|������������� ��50BT}x ������ ,UPbt�� �����/-/(/ :/L/u/p/�/�/�/�/ �/�/? ??$?M?H? Z?l?�?�?�?�?�?�? �?�?%O O2ODOmOhO zO�O�O�O�O�O�O�O 
__E_@_R_d_�_�_|�_%�C_RPI<�N�_�_"oo�_;���_.owo�o�o(�SL�_@l`�o�c�o  $;HZl��� ������ �2� D�[�h�z������� ԏ���
��3�@�R� d�{�������ßП� ����*�<�S�`�r� ��������̯��� �+�8�J�\�s����� ����ȿڿ���"� 4�K�X�j�|ϓϠϲ� �o�fYo�a�o�o�+� =�O�a�s߅ߗߩ߻� ��������'�9�K� ]�o��������� �����#�5�G�Y�k� }��������������� 1CUgy� ������	 -?Qcu��� ����//)/;/ M/_/q/�/�/�/�/�/��/�XNOCODE� H]e��GkPRE_CH�K J]k� A �� �< ��� ]ee?w?]e 	 <Y?�?�?�Ù?�? �?�?O+OOOaOsO MO�O�O�O�O�O�O�O _'__K_]_7_�_�_ �?{_�_�_u_�_o�_ oGo!o3o}o�oio�o �o�o�o�o�o�o1C gyS���_�_ ����-���c� u�O���������ᏻ� ͏�)��M�_�9�k� ��o���˟ݟ���� ���I�[�5����k� ��ǯ��������3� E��i�{�U�g���ÿ �����ӿ�/�%�� e�w�ϛϭχϹ��� �����+��O�a�;� mߗ�q߃����߹�� ���!�K�A�Sρ�� -����������� 5�G�!�S�}�W�i��� ����������1 gyS��i� ���-Qc =O������ //�/M/_/9/�/ �/o/�/�/��/?? �/7?I?#?U??Y?k? �?�?�?�?�?�?	O3O OOiO{OUO�O�O�O �O�O�/�/_/_�O;_ e_?_Q_�_�_�_�_�_ �_�_o�_oOoao;o �o�oqo�o�o�o�o �o9K_3�� m������� 5�G�!�k�}�W����� �������Տ�1�� U�g�]O�����I�ӟ 埿������Q�c� =�����s���ϯ���� ���;�M�'�Y��� y�����˿e�׿�ۿ �7�I�#�m��Yϋ� �Ϗϡ�������!�3� �?�i�C�Uߟ߱ߋ� ���ߡ����/�	�S� e�?���u������ ������=�O�)�;� ����q��������� ����9K��o�[ �������# 5AkEW�� �����/' U/g//s/�/w/�/�/ �/�/	??�/'?Q?+? =?�?�?s?�?�?�?�? O�?�?;OMO'OqO�O =/kO�O�O�O�O_�O %_7__#_m__Y_�_ �_�_�_�_�_�_!o3o oWoioCo�o�o�O�o �o�o�o�o)S -?��u��� ����=�O�)�s� ��_������o�o�� ���9��%�o���[� ������ß�ǟٟ#� 5��Y�k�E�w���{� ��ׯ�ï��ُ� U�g�A�����w���ӿ ����	����?�Q�+� uχ�a�sϽ��ϩ��� ���)�;�1�#�q߃� ߧ߹ߓ��������� %�7��[�m�G�y�� }���������!��� -�W�M�_ߍ���9��� ��������AS -_�cu��� ��=)s �_��u���/ �'/9//]/o/I/[/ �/�/�/�/�/�/?#? �/?Y?k?E?�?�?{? �?�?��?OO�?CO UO/OaO�OeOwO�O�O �O�O	_�O_?__+_ u_�_a_�_�_�_�_�_ �?�?)o;o�_GoqoKo ]o�o�o�o�o�o�o�o %�o[mG���}�����!�����$DCS_S_GN KeM���w@5a0�7-NOV-20 00:43 ��10-JUL�-18 22:4�9g����� Q=�����������R�S]���Z�o��5�ڞ� � 9�VERSIO�N E�V�4.2.10ϋE�FLOGIC 1�Le�  	���`)��`8��PROG_�ENB  ��� ���Y�ULSE � >�q��_A�CCLIM����s����WRS�TJNT��M��5�EMOb���u�
��ݐINIT M��jזOPT_�SL ?	f�
� 	R575���C�74H�6I�7RI�5��s�1m�2I��*����&�TO  �2�����V��DKEX��dM���(�PATH AE��A\ D\  ?\ \IMGB�M��_���HCP_CL?NTID ?� � *�����؂�IAG_GRP �2Re� ���`E��  F?h F�x E?`��D�����B�  �Ϣ����A�/�C�f  Cyj�Y��dCj�q�B��i���mp�3m6 7890?123456����`�  A��ffA�=qA��  AхAʯ�HAľ���������A���������@���g�A�p�����A����g�B4�� 袅2���
���(��A�A�
=�A�B���A���
A�Q�A�:�������j������j!�	n5��W{A�Z�̶��Z����������A�:��������h�z���ߞ߰�6�EG�A}@��:�RA5Z�U/��)��#F�Z�b�������*�<�>6�Pz�AJ��Y��?��9p�A3\)A,��A&����~�������4�cF�]��AW���P��J��C��<�Z�4��-Z�%G� ��0�B�T�6�%�
 	n��?Q��%o� w��Yk�)@M_�kc���Q���i�����=׿
==�G��>�Ĝ��7'�=��6�7����@ʏ\&�p�4$%��@�Ah��/ �A��<i��<�xn;=R�=�s��=x<�=��~Z�;��|%<'�'������?+ƨC�  �<(�U�� 4�"����&����%��\က?ň? �?6?H?h�$T?~?�?�?�?�?�?�?�?)7L?S�FB'$�/Eͽ�4OG�ΐ
Ա��iDj�L�x�CA��G�X�j�|�챤��O�L����Oʹ�%_sNED�  E�  Eh'� DQPXR:_�� �_���u�_�_�_��q_�_m_o�K4o:b���D�|-�0���C3u|����À�B�T�o�o o�o�o�o�o��o��E}�?��"� _r>���>im����Y<�=<��Du;ě�Pu��C�T_CONFIG� S׷񓄄�eg?�ʱST�BF_TTS��
@q��s�������v9��MAU��f�x�MS�W_CFtpT׻ � ΌOCVIE�W�pU���� �_Y�k�}��������r G�܏� ��$�6�ŏ Z�l�~�������C�؟ ���� �2�D�ӟh� z�������¯Q���� 
��.�@�ϯd�v��� ������п_����� *�<�N�ݿrτϖϨ�X����\|RC �V�5�r!h��^�9�(�]��L߁�pߥ��tSBL�_FAULT �W�����GPMSqK�w��hpTBR �#X��>��q�o�xF�X���TDIA	�Yxy��sM!�UD1: 6�78901234!5��rM!��P(��� ��	��-�?�Q�c�u� ���������������F��	�"
��Mt�ORECP���
�� ��������  $6HZl~�� ����#52/���UMP_OPTGION�p��R!T�t�s��s%PME�u�f/Y_TEMP � È�3B�̈p� �A� �$UN�I�p�u�!��YN_?BRK Z2��?EDITORX!^!��/2_j ENT �1[��&�,&�JR_SETUP�PROGRAM 9H�pmpHEC����&HOME J�ACKPO:0IG�h?�u&MAI�N�?�? &P�ICK_�?�?#&�:LEF�p�?���&PNS000�1 OSE E ��?x8CLAV C�L<Or<&GRIPPE�gBnO��&X0CALI'CRA["] T�O�C�CAMEA�BB8�D�O�r&�H�C��@�O�p&PLGACE�<$_�p_�0�=ZBHP_�pd&�X1HIP FTH�BE�A}_1W4A�_�t=ZERO 9@PALLET_H�_�z6<PSTIC_��_�\/&CLE?AR_IO �F�p��4t<gT dYeYo�&�	MID_POI�@0$`B�Ѕo  �0MGDI_ST�A�%<q�! � m+0NC�c1\�� ��"~
"~d(/o���� �����#�5�G� Y�k�}�������ŏ׏ 鏀% ��$�6�D�\q D�j�|�������ğ֟ �����0�B�T�f� x���������үL��� ��'�9�S�]�o��� ������ɿۿ���� #�5�G�Y�k�}Ϗϡ� �����������1� K�U�g�yߋߝ߯��� ������	��-�?�Q� c�u��������� ����)�C�9�_�q� �������������� %7I[m� ��������! �M�Wi{��� ����////A/ S/e/w/�/�/�/�/� ��/??+?EO?a? s?�?�?�?�?�?�?�? OO'O9OKO]OoO�O �O�O�O�O�/�O�O_ #_=?G_Y_k_}_�_�_ �_�_�_�_�_oo1o CoUogoyo�o�o�o�o �O�o�o	5_'Q cu������ ���)�;�M�_�q� ���������oŏ�� �-?I�[�m���� ����ǟٟ����!� 3�E�W�i�{������� ˏݏ�����7�A� S�e�w���������ѿ �����+�=�O�a� sυϗϩ�#�կ���� ��/�9�K�]�o߁� �ߥ߷���������� #�5�G�Y�k�}��� �����������'�1� C�U�g�y��������� ������	-?Q cu������ ��;M_q �������/ /%/7/I/[/m//�/ �/���/�/�/�/) 3?E?W?i?{?�?�?�? �?�?�?�?OO/OAO SOeOwO�O�O�/�/�O �O�O_!?+_=_O_a_ s_�_�_�_�_�_�_�_ oo'o9oKo]ooo�o �o�o�O�o�o�o�o_ #5GYk}�� �������1� C�U�g�y������o�� ӏ����-�?�Q� c�u���������ϟ� ���)�;�M�_�q� ��������˯ݯ�	� �%�7�I�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϧ��� ����������/�A� S�e�w߉ߛ߭߿��� ������+�=�O�a� s���ϱϻ������� ��'�9�K�]�o��� �������������� #5GYk}��� �����1 CUgy���� ���	//-/?/Q/ c/u/�/��/�/�/�/ ��/?)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�/ �/�O�O�O�O?_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_oo/oAo Soeowo�O�O�o�o�o �o�O+=Oa s������� ��'�9�K�]�o��� �o����ɏۏ�o��� #�5�G�Y�k�}����� ��şן�����1� C�U�g�y��������� ӯ�߯	��-�?�Q� c�u���������Ͽ� ���)�;�M�_�q� ��}ϧϹ������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�ϕϟ�� ����������/�A� S�e�w����������� ����+=Oa ��������� '9K]o� �������/ #/5/G/Y/k/��/�/ �/�/��/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cO}/kO�O�O�O�/�O �O__)_;_M___q_ �_�_�_�_�_�_�_o�o%o7oIo[ouO ��$ENETMOD�E 1]�E��  �@��@�a�D�o�`|hR�ROR_PROG %�j%F�oy��eTABLE  �k�OCUguw��bSEV_NUM� �b  ���a�p�a_AUT�O_ENB  ��e�c�d_NO�q �^�k�a�r W *��p��p��p	��p�p+�p��,���tFLTR��vH�IS�s�A�`�{_A�LM 1_�k e��D�|@+-��ȏڏ����"�1�_\�r�p  �k�q��bg��`TCP_V_ER !�j!�o�2�$EXTLOGo_REQh��yι�SIZ��ST�Kߙ�u���T�OL  �ADz�p��A ��_BWDG��L�H��b1��DI6� `�E�L��d�AM�ST�EP^�p��`��OP�_DO��aFAC�TORY_TUN�h�dɩDR_GR�P 1a�iR�d �	b� ��`��������gl�rw�q�����J ���T��f�w�a����� �����Ϳ���<�x'�`�K�<��>�E�<`~�=�īf
 Ifٓ�Ϲ�`��C��������	�C`�}dC��N<�B��{D� �@UU�T`�UT ߉�$� _E�� �߀���OHcEP]���O��#M��^��KA��x�?��� ��:6:N{�,�9-�4��x�
( ���� m-���!o���b�e�3�
{FEATURE� b�EH��a�HandlingTool ����BEngli�sh Dicti�onary��4Dw St��ard�����Analog �I/O����gle� Shift��u�to Softw�are Upda�te�matic Backup���E�ground �Edit���Ca�mera��F��CnrRndImJ����ommon calib UI|���nc��Moni�tor��tr��R�eliab��D�HCP����ata Acquis��~��iagnosA����ocument Viewe�����ual Che�ck Safet�y���hance�d����s` Fr�t��xt. DI�O ��fiD�e�nd� Err��L(C��s�	r��� � 7���FCTN /Menuy v��*�TP Infayc@��GigER�d\�p Mask� Exc� g�H�TPProxy �Sva�igh-wSpe� Ski����< � mmuni�c@�ons�ur�7	��Scon�nect 2	(n{crRstru��$*0 eWq JC���KAREL Cmod. L�ua�~g#Run-Ti� �Env](el u+D�sB�S/W��Licenses�`� Book(S�ystem)��M�ACROs,�/�Offse��%H0� *�� MR�����BMechStoEp�t  (�%i��	�\6x� ��B�>o}d�witch�?�037.6�;Optqm�?03�fil`�/7g��%ulti�-T�f��PCMO fun:'8Io%xt1DXMRegi� Yr�;FriY FHK��F��Num Se�lT5�I�  Adj�u��N�A	��Mta�tu�A�O[
��RDM Robot���scove��8Ue�a)@� Freq �Anly�Rem�R0�n��8UDRSe�rvo� �0��SN�PX b�"�SN�PCliX�^
�LGibr���_�� c4��P�Vo� t7ss#ag1E��{� �1̡�{�/IQ4eMI�LIB]o7bP F�irm(�GnP7A�cc]�e�TPTX5deln0zo8ax�� 5Hmorqu�imula��z��fu�0Pa�!Gn\���:�3&�ev.4e ��riq �oUSB� port ��i�P� aY �vR E�VNTw�pnexcept� yPfD�u,��VC��r��X8V$ ��o��[��S�PSC�eH�SG�E]�S�UI��Web PlV���Q�ང��WZDT Appl���v����GridHQp�lay�D`I�&�R��r.��`�7�;R-�2000iC/1�25L��2D G�ui�pZ����Gr�aphic����D�V- Path Ctr��������dv�DCS<pc�kw!��larm �Cause/wPe}d��Ascii���BLoad` \�Usplr��toS���%prityAvo�idM��l����GAu�氯¢8���s��t����yc��"�@�rp~ ��5�os./�cu �z��%	�trans.be�tw.CRLmai�n N��Q.��t?herNetZaz���`��ca ��,RA<p� ��(&0~Q/C�@o�'���L�<�o�89���NRT쫖�On��e H�el��<E�@�AQ�t=r�ROS ��7��e퇟� ����s�up�rt���vH�apA�[����Pk��GiG� t�݋Im�0F�0X�P�n�sp !+�|�64M?B DRAMdώӇFRO�����l�e3ll���sh����"�c�;��%�p>v�ty�s�B��� r �B��_R�0���~Ѐ3���hxP���MAIL⋞}�r �[ЄCP�R��q�T1���[��!Adp.G�X�s����/4Lz�arHQq�Z�%�Ro��+ax���OGPT Pؿ�Ac'`���TX!qpXpSyn�.(RSS)TVquir<`��DR�UpT��^� (�uess��S���]�V�RS6�dauXp�[?��Pmi��3DLb�^�w!�e��K�`l Bu�i)@n�APLCdKV�Հ�CGUNxCRG���DD@̪�LS���BU����K�! /V�TA�T*&B��C*^�X/TCBm/&4/~'x�~'F�/&p~'�
7�u?TEH1?C6�B7!Vi?C6\�
6FP/�7l/
6G�/�7�?�7?2
6H,O
6IAIO[FLHO
6LN�O+%MO �G�/�G/
6N�O
6!PdOW�?
6R�?
6!SD_rW`_
6W�_�W�_
4VGF�_�UP�2��W�O�W�_�VB$@o�VD\o�VF�/�V�O�TUT<b01�o�f2�o�bTBG�G$b�lr~��� U9I�`|�HMI"r��pon��`�Q�fo�r s�>s�KARcELK��al�TPY��c|��|����� �����*�<�i� `�r�������Տ̏ޏ ���&�8�e�\�n� ������џȟڟ��� �"�4�a�X�j����� ��ͯį֯����� 0�]�T�f�������ɿ ��ҿ������,�Y� P�bϏφϘ��ϼ��� ������(�U�L�^� �߂ߔ��߸�������  ��$�Q�H�Z��~� �������������  �M�D�V���z����� ����������
I @Rv���� ���E<N {r������ �//A/8/J/w/n/ �/�/�/�/�/�/�/�/ ?=?4?F?s?j?|?�? �?�?�?�?�?�?O9O 0OBOoOfOxO�O�O�O �O�O�O�O_5_,_>_ k_b_t_�_�_�_�_�_ �_�_o1o(o:ogo^o po�o�o�o�o�o�o�o  -$6cZl� �������)�  �2�_�V�h������� ˏԏ���%��.� [�R�d�������ǟ�� П���!��*�W�N� `�������ï��̯ޯ ���&�S�J�\��� ��������ȿڿ�� �"�O�F�Xυ�|ώ� �ϲ���������� K�B�T߁�xߊ߷߮� ���������G�>� P�}�t������� �����C�:�L�y� p�������������	  ?6Hul~ ������ ;2Dqhz�� ���/�
/7/./ @/m/d/v/�/�/�/�/ �/�/�/?3?*?<?i? `?r?�?�?�?�?�?�? �?O/O&O8OeO\OnO �O�O�O�O�O�O�O�O +_"_4_a_X_j_�_�_ �_�_�_�_�_�_'oo�0o]oTol  ?H552oc�a�21�eR78�h5�0�eJ614�eAwTUP�f545�h�6�eVCAM�eC�RI�gUIF�g2�8�fNRE�f52��fR63�gSCHޛeDOCVOvCS]U�f869�g0�f�EIOC+w4�fR{69�fESET�gv�gJ7�gR68�f�MASK�ePRXuYx7�fOCO�x�3�h�f�p�h3�vJ�6�h53rvH$�L{CH�vOPLG�g�0�MHCR�vS�m�MCS�h0�w5=5�fMDSW���;OP�MPR�?p�2�0�fPCMvR�0���p�fw�2�51��g51.�0�fPR�S�w69�vFRD��fFREQ�fMC�N�f93�fSNByA7w%�SHLB���M��?p��2�fHT=C�fTMIL�hrv�TPA�vTPTXF�EL��w�rw8�gܯ`�fJ95vTU�T�95�vUEV�vUEC�vUFR��fVCC��O��V�IP��CSC�C�SG*vdpI�eWE�B�fHTT�fR6l5x@�CG��IGݧoIPGS�RC���DG�H72�w9nQ�R76�fR8���w�b�85rvR66tb��wR,�R51�w�53"�68n�66��2�6.�6vJ74�g75b���`�b�<�R5Y�J59�.�58.�85�54���6m�NVD�vR�6y����87j�40v�p:�i�R7w�p�vD0m�F�RT�S��CLI��gC�MS�v?��fSTY:��6��CTO�fcpڊw7qxNN
�NN��vORS���pF�3:��5�HPM�z�8\�?p�fOPI2�3кڸ7rvCPR��LꡧS��7�vSVS�NvSLM�vV3Dܺ�wPBV�AP�L�vAPV�CC�G�fCCRn�CDCDL2�CSBnfvCSKCT��CTBަ�TCh�����CҧTCvl��TC��TC�v�CTENvs��TEXZvs�ƧTF
�F��G��G��^�H^�I��T�CT)�CT�M��� ��N^�P���P��R
�A�TSr
�Wr	2�VGF�P2��P2��� �UB�D�FvV��VT�g� �fVTBZ��VewIH�V;�
K��V��vhQc u������� //)/;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m??�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S��e�w�  H55y�����R78��50��Jw614��ATU�����545��6��VsCA���CRI��UI���28�N�RE��52�R6�3��SCH��DO�CV��C��86u9��0��EIO2�e�4��R69�EgSET���J7��R68��MASK^��PRXY?�7��OCO3��� ���3n
J6��53���H�LCHN
O�PLG��0�
MH�CRO
SMCS���055��MD�SWo}OP}M�PR~
{�0��PCM>�R0� ��l�51��51,�0��PRS69�n
FRD.�FRE�Q��MCN��93���SNBAo��SHLB�*M�+{�^�2��HTC��TMsIL���TPA��oTPTX:EL�*���8���~�J9�5N�TUT~95�n
UEV
UEC�N
UFR.�VCC��<O.VIP:C;SCN:CSG^����I��WEB��HT�T��R6m�|<CG�mKIGMKIPGS��JRC:DG}H�72��9=+R76���R8]P�K85N��R66�L��R,�R51��53�6�8[66�2�6�,6N�J74��7�5�L����K�R5n�;J59k58k�8m<54n[6[NVD
R6[P�87^l4N�; l]+cR7M�; N�D0[�F,|RTS�*CL9I���CMS��{p���STY;6mC�TO�����7��N�N�[NNn
ORS�.; .l3�k5�[H�PM�L,{���O�PI�Jkp�\7��C�PR~+L�;S�7�n
SVS��SLM�
V3DL=�PB�VN:APL��AP�V~
CCG��CC�RCD�;CDL�JCSB��CSKv~CT=;CTBNJ�ېKTC�*��ΜC�>KTC>���^�TCv��TC
CTE���k�n�TE��k�.KTUFޜF�GΜG���N�HN�IN{T��CT];CTM�M�;����NN�P�PΜR,ޜ}|TSޜW���J�VGF޻P2�;PQ2�*���B�D�5F>�V��VT��k����VTB~�V��I�H;V�@��KKV mJ~�����	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q����������� ��%�7�I�[�m�� �������������� !3EWi{�� �����/ ASew���� ���//+/=/O/ a/s/�/�/�/�/�/�/ �/??'?9?K?]?o? �?�?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_ �_�_�_�_	oo-o?o Qocouo�o�o�o�o�o �o�o);M_ q������� ��%�7�I�[�m�� ������Ǐُ���� !�3�E�W�i�{����� ��ß՟�����/� A�S�e�w��������� ѯ�����+�=�O� a�s���������Ϳ߿ ���'�9�K�]�o� �ϓϥϷ��������� �#�5�G�Y�k�}ߏ� �߳�����������1�C�U�g�y����STD��LANG�������� �����"�4�F�X�j� |��������������� 0BTfx� ������ ,>Pbt��� ����//(/:/ L/^/p/�/�/�/�/�/��/�/ ??$?6?H4R{BT��OPTN_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO��O�O�O�O�O�ODPN��	__-_?_ Q_c_u_�_�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m �������� !�3�E�W�i�{����� ��ÏՏ�����/� A�z�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo�%o7oIo[omod9�9{e�$FEAT�_ADD ?	�����a�`  	zh�o�o�o �o'9K]o �������� �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� ��ӟ���	��-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������� #5GYk}� ������// 1/C/U/g/y/�/�/�dDEMO b�i?   zh�- �/�/??"?O?F?X? �?|?�?�?�?�?�?�? OOOKOBOTO�OxO �O�O�O�O�O�O__ _G_>_P_}_t_�_�_ �_�_�_�_oooCo :oLoyopo�o�o�o�o �o�o	 ?6H ul~����� ���;�2�D�q�h� z�����ˏԏ��� 
�7�.�@�m�d�v��� ��ǟ��П�����3� *�<�i�`�r�����ï ��̯����/�&�8� e�\�n���������ȿ �����+�"�4�a�X� jτώϻϲ������� ��'��0�]�T�f߀� �߷߮���������#� �,�Y�P�b�|��� �����������(� U�L�^�x��������� ������$QH Zt~����� � MDVp z������/ 
//I/@/R/l/v/�/ �/�/�/�/�/??? E?<?N?h?r?�?�?�? �?�?�?OOOAO8O JOdOnO�O�O�O�O�O �O_�O_=_4_F_`_ j_�_�_�_�_�_�_o �_o9o0oBo\ofo�o �o�o�o�o�o�o�o 5,>Xb��� ������1�(� :�T�^����������� ʏ��� �-�$�6�P� Z���~�������Ɵ� ���)� �2�L�V��� z�������¯���� %��.�H�R��v��� ����������!�� *�D�N�{�rτϱϨ� ����������&�@� J�w�n߀߭ߤ߶��� ������"�<�F�s� j�|���������� ���8�B�o�f�x� ������������ 4>kbt�� ����0 :g^p���� ��	/ //,/6/c/ Z/l/�/�/�/�/�/�/ ?�/?(?2?_?V?h? �?�?�?�?�?�?O�? 
O$O.O[OROdO�O�O �O�O�O�O�O�O_ _ *_W_N_`_�_�_�_�_ �_�_�_�_oo&oSo Jo\o�o�o�o�o�o�o �o�o�o"OFX �|������ ���K�B�T���x� ������������� �G�>�P�}�t����� ����������C� :�L�y�p��������� �ܯ���?�6�H� u�l�~��������ؿ ���;�2�D�q�h� zϧϞϰ������� � 
�7�.�@�m�d�vߣ� �߬����������3� *�<�i�`�r���� ���������/�&�8� e�\�n����������� ������+"4aX j������� �'0]Tf� �������#/ /,/Y/P/b/�/�/�/ �/�/�/�/�/??(? U?L?^?�?�?�?�?�? �?�?�?OO$OQOHO ZO�O~O�O�O�O�O�O �O__ _M_D_V_�_ z_�_�_�_�_�_�_o 
ooIo@oRoovo�o �o�o�o�o�o E<N{r��� ������A�8� J�w�n���������Џ ڏ����=�4�F�s� j�|�������̟֟� ���9�0�B�o�f�x������ȭ   ��ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6HZ l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/�l/~/�/�/�/�)  �(�!�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>Pbt� �������� (�:�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτϖ� �Ϻ���������&� 8�J�\�n߀ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x��������������� ,>Pbt� ������ (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?V? h?z?�?�?�?�?�?�? �?
OO.O@OROdOvO �O�O�O�O�O�O�O_ _*_<_N_`_r_�_�_ �_�_�_�_�_oo&o 8oJo\ono�o�o�o�o �o�o�o�o"4F Xj|����� ����0�B�T�f� x���������ҏ��� ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ ؿ���� �2�D�V� h�zόϞϰ������� ��
��.�@�R�d�v� �ߚ߬߾�������� �*�<�N�`�r��� �����������&� 8�J�\�n��������� ��������"4F Xj|����� ��0BTf x������� //,/>/P/b/t/�/P�/�/�/�!� �( �/�/
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�o�o �o�o�o0BT fx������ ���,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� �ߨߺ��������� &�8�J�\�n���� �����������"�4� F�X�j�|��������� ������0BT fx������ �,>Pbt �������/ /(/:/L/^/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n��� ������"�4� F�X�j�|�������ď ֏�����0�B�T� f�x���������ҟ� ����,�>�P�b�t����������Ω�$F�EAT_DEMO�IN  Ӥ�����Ԡ�IND�EX����I�LECOMP �c���4����*�SETU�P2 d4�~>��  N i��'�_AP2BCK� 1e4�  #�)Ϩ����%��пԠ7�����ѥ��'� ��K�ڿXρ�ϥ�4� ����j��ώ�#�5��� Y���}ߏ�߳�B��� f�����1���U�g� �ߋ�����P���t� 	����?���c���p� ��(���L������� ��;M��q �� 6�Z�~�%� I�m�2� �h��!/3/�W/ �{/
/�/�/@/�/d/ �/?�//?�/S?e?�/ �??�?�?N?�?r?O �?O=O�?aO�?�O�O &O�OJO�O�O�O_�O 9_K_�Oo_�O�_"_�_��_C�w�P{� 2>��*.VR�_o�P*oCo�SIomo�WU`PCuo�o�POFR6:�o�nYo�o}kT�$�e�N|���otVV*.Fo��Q	�c��|qa��{STM� +��b�`�V��z��{HG���<���X�j����zGIF	�3�>���܏��zJPG ����>���`�r��~j#JS�:��P͓(���%
JavaS�criptf���C�SW���=���h� %�Cascadi�ng Style Sheets��\P
ARGNAMOE.DT�|\A��\-��M�]�n��>]�DISP*d�G��A���񿀵�򿞿
�TPEINS.X3ML!�Ϳ:\5���U�Custom Toolbarv����PASSWOR�D�z^FRS:�\��x� %Pa�ssword Config�Ϧ����Y�@���ϥ�W_ ��{_���߱_#��G� Y���}����B��� f������1���U��� y������>�����t� 	��-?��c��� ��L�p �;�_q �$ ��Z�~/�/ I/�m/��/�/2/�/ V/�/�/�/!?�/E?W? �/{?
?�?.?�?�?d? �?�?O/O�?SO�?wO �OO�O<O�O�OrO_ �O+_�O$_a_�O�__ �_�_J_�_n_oo�_ 9o�_]ooo�_�o"o�o Fo�o�o|o�o5G �ok�o��0�T �����C��<� y����,���ӏb��� ���-���Q���u��� ���:�ϟ^�ȟ��� )���M�_����� ��H�ݯl�����7� Ư[��T��� ���D� ٿ�z�Ϟ�3�E�Կ i����ϟ�.���R��� v���߬�A���e�w� ߛ�*߿���`��߄� �+��O���s��l� ��8���\������'� ��K�]���������� �$FILE_�DGBCK 1e�������� < �)�
SUMMARY�.DG��e�MD�:��-q�Di�ag Summa�ry.;�
CONSLOG#q��@Conso?le log�:�	TPACCN��%�1<TP� Account�in�;�FR6�:IPKDMP.'ZIPei�
}��=MExcept�ion�;�*.�DT�/q�FR�:\�>.�FR� DT File�s>/j MEMCHECK'��/��Memory� Data�/���(i\)�!RIP�E��/�/A?�#%�1 Packe�t L��%�b<"1STAT;?"?|4?�? %]2�Statu_/y<	FTP?!O�?%O�'��mment �TBDNO�'���)ETHERN�E�?&O�!�O�O@?Ethernf0� ?figura�A�~8ADCSVRFBO�(O:OS_�3P v�erify al�lV_�$���UDIFFK_1_C_�_W3mXdiff�_�W�!>PCHG01�_�_��_]o�1�_�o�R�i2So:oLo�o�_�o��o"b3�o�o�oe� �o�vVT�RNDIAG.LAS�BT��!�qO Ope�Ch1 E�nostic�'���<)VDEV�rDA0/��m��1�Vis�Dev�ice� �IMG@�r�H�Z��V3���Imag���U�P6�ES5�ʏF�RS:\5�@/B U�pdates L�istv�;�݀FLEXEVEN�O�Ώ�����1�� UIF EviAi?�#��Ѱ)
PSRBWLD.CM%��e�a�=�x�� PS�_ROBOWELoO9��AIOׯ�����'�BNet/�IP�pa"��#ߌ�)�GRAP?HICS4D������%4D �Graphics�Z/�'�' 2GI�G?�o���&G�igE���#���2SMOc�����'P�/Emai�l$�=��\��SHADOW��h�z����#Shadow? Chang���&� ﾣRCMERAR����ϓ��#X��CFG Erro�r��t��6� ��+��3CMSGLIB��r߄�������2�������*�)�ZDT�s���n�'ZD0�ad9����&쿢NOTI�_v����%Notific�B���&�A�)��u�X�d��������������� ������AS��w �*<�`� �+�O�H� �8��n/�'/ ��]/��/�/"/�/ F/�/j/�/?�/5?�/ Y?k?�/�??�?B?T? �?x?OO�?CO�?gO �?`O�O,O�OPO�O�O �O_�O?_�O�Ou__ �_�_:_�_^_�_�_�_ )o�_Mo�_qo�oo�o 6o�oZolo�o%7 �o[�ox�D �h���3��W� �������ÏR�� v�����A�Џe�� ����*���N��r��� ���=�O�ޟs���� &���ͯ\�񯀯�'� ��K�گo������4� ɿۿj�����#ϲ�� Y��}�ϡϳ�B��� f��ϊϜ�1���U�g� �ϋ�߯�>ߨ���t� 	��-�?���c��߇���(��x��$FI�LE_FRSPRT  ����������MDONLY 1�e��|� 
 ��)MD:_V�DAEXTP.Z�ZZ��z�Q�`��6%NO Ba�ck file <+�B��U�W�� A�������Q�0�� Tf�����O �s�>�b �o�'�K�� �/�:/L/�p/� �/�/5/�/Y/�/}/�/ $?�/H?�/l?~??�? 1?�?�?g?�?�? O2O~��VISBCK	�|���*.VD3O|}O�0FR:\L@�ION\DATA�\hO�2�0Vision VD~���O�8*.CAM�O_ %	�A�C�O��LGigE C�amera Definit�@-_�? }_�?�_O�_�_f_�_ �_o1o�_Uo�_yo�o o�o>o�o�oto	�o -�o&c�o�� �L�p���;� �_�q� ���$���H� ���~����$�I�؏�m�7NLUI_CONFIG f���_A|� $ 	Z��{��ӟ���`	��-�;���|xc� e�w���������S�� ���(���9�^�p� ������=�ʿܿ� � �$ϻ�H�Z�l�~ϐ� ��9���������� � ��D�V�h�zߌߞ�5� ��������
���@� R�d�v���1���� ��������<�N�`� r�������������� ��&8J\n� ������� "4FXj|� ������/0/ B/T/f/x//�/�/�/ �/�/�/�/?,?>?P? b?t??�?�?�?�?�? w?�?O(O:OLO^O�? �O�O�O�O�O�OsO _ _$_6_H_Z_�O~_�_ �_�_�_�_o_�_o o 2oDoVo�_zo�o�o�o �o�oko�o
.@ R�ov����� g���*�<��M� r���������Q�ޏ�� ��&�8�Ϗ\�n��� ������M�ڟ���� "�4�˟X�j�|����� ��I�֯�����0� ǯT�f�x�������A��Robot S�peed 10%��������1�?��H�x8�E��$FL�UI_DATA �g���u��?�g�RESULT 2hu���� �T��/wizard�/guided/�steps/ExpertT������� ��/�A�S�e�w߉�����Skip �G��ance a�nd Finish Setup�� �������"�4�F�X�pj�|��<� H��.?�uŷ�0� �H�����u����ps��"�4�F�X� j�|������������� ��H�!3EWi {������?�@��?�����+��&���rip����Too�lNum/NewFrame��� �����//*/<</��0x0?/g/ y/�/�/�/�/�/�/�/p	??-???  <��;?����di�meUS/DST B?�?�?�?OO/OAO�SOeOwO�O��Enablv�O�O�O�O __)_;_M___q_�_
�_F�G��?q?�_�?�?�224�?%o7o Io[omoo�o�o�o�o �o�O�O!3EW i{��������_�_�_,��_ ozon�0�}�������ŏ�׏�����1����EST Ea��rn St�Э�;�t� ��������Ο����`�(�:���J� �?��7��{���Ϻ�Region>�ͯ߯ ���'�9�K�]�o������America���Ϳ߿�� �'�9�K�]�oρ�@�R�y�i����ϟ�b?Editor��!� 3�E�W�i�{ߍߟ߱����������ula�r 
�� (re�commen�) ��(�:�L�^�p��� �������G��������#�����/acces��t����������������(?��Connect �to Network7n���� ����"4K�a����s��!I��_�Introduct�����// &/8/J/\/n/�/C�p �/�/�/�/�/�/?? 0?B?T?f?x?�?�rR���r�i�?9��/Safet��O O2O DOVOhOzO�O�O�O�O �O�/�O
__._@_R_ d_v_�_�_�_�_�_�_ �?�?�_'o�?W�j�oo �o�o�o�o�o�o�o�o #�OGYk}� ��������@1��_oov�8i#Eo�Wf/current8�͏ߏ���'��9�K�]�o���D15�-MAY-20 �09:31 AM ����П�����*�@<�N�`�r������球�e�ǯ5l ����Yea��/�A�S�e��w���������ѿ@2020ۿ��(� :�L�^�pςϔϦϸ������ 
����  �䷯ߋ��Month��s߅ߗ� �߻���������'�B5/�U�g�y�� �����������	��-����� �m�3nA߫�DaO���� ����0BTfx��1C��� ��'9K]o�@�R�_��ۯ����Hou�/+/ =/O/a/s/�/�/�/�/�/8�9�/�/?!?3? E?W?i?{?�?�?�?�?��?�R�	�O3n"|�S�inute�? pO�O�O�O�O�O�O�O0 __$_�31+_R_ d_v_�_�_�_�_�_�_@�_oo*o�?S�Opio�=O��AMP�� �o�o�o�o	-? Qcu������ ����"�4�F�X��j�|�����攠�{o]o��-L�o��NetDon^O�#� 5�G�Y�k�}������� ş�Z������1� C�U�g�y���������ӯ8aCo����;��&�ripper�O�oolNum/FraX�s �o��� ������ɿۿ���� #�>�@_L�^�pςϔ� �ϸ������� ��$�@;oQ����i�/J)9�~K�ActiveW� *����������!�3��E�W�i�(�0x0 {�������������!�3�E�W�i�{�  �=��������ߗ�MOacroS���w��s~�-?Qcu ����|��� );M_q�� ���������/.K�,������Open \�o/�/�/�/�/�/�/ �/�/?�:�G?Y?k? }?�?�?�?�?�?�?�? OO6�H�/dO֏�Summary&O �O�O�O�O�O_"_4_ F_X_j_ٟ�_�_�_�_ �_�_�_oo0oBoTo foxo��[O�oO�RobotOp|o 
.@Rdv� ���}_���� *�<�N�`�r����������̏�o�o�o��f-|5/G/oClos[� k�}�������şן�����2�E�W� i�{�������ïկ� ����4OFI��]���n1��BetMethod"���ǿٿ ����!�3�E�W�i��,7Direct� entry o�f EOAT datasϱ������� ����/�A�S�e�v��]�RB�U����h�$���Btraig�htOffset v�� �2�D�V�h�z�����12�� Tool������ /�A�S�e�w����������~���ߤ��m%�ߚA��AX��cu ��������21298.4993�GYk}� ������/-y5�C�?���]/1CY/�/�/ �/�/�/?#?5?G?Y?�k?�q	-169.1565o?�?�?�? �?�?�?	OO-O?OQO�cO"/4/���)( O/�Os/�/CZrO_ _/_A_S_e_w_�_�_��_�_*951.8884�_�_oo&o 8oJo\ono�o�o�o�oxuO�O�CDm�ۣO���)�O��Rot_ation=wW�o cu����������_179.868�?C�U�g�y� ��������ӏ���	�8�o�oD%3�V�oY�-?P���ɟ۟ ����#�5�G�Y��-.2586k� ������̯ޯ����&�8�J�\��-�g���hK���o�����Rn���/�A�S�e��wωϛϭ�l�-2?9.4700���� ���"�4�F�X�j�|���ߠ߲�q�������#����J"ѿ��tp3Zdir/Tp3z��X�j�|� ������������� �_0�B�T�f�x����� �������������ߐ�o�_Ͱ+%��M�easureme�nt/Straigh�O����� 1CU�&�� ������	// -/?/Q/c/"4F�/�j|/We�Nu�ms/New�#s j/	??-???Q?c?u?p�?�?�?j0x�� �?�?OO*O<ONO`O@rO�O�O�O�Op}/��I�/�O�.�/�,Twool�#Use�O `_r_�_�_�_�_�_�_�_om1o5oGo Yoko}o�o�o�o�o�o�o�op
�OQp��OM_!_�,PartF_��������)�;�M�_�b2 c���������я��� ��+�=�O�a� 2y�?���(u�'s/Gڰ�#f���&� 8�J�\�n����������71.10�� ����)�;�M�_��q���������|/�&BG�33�����)ɟ�ۙPayload1Cm�V�h�zόπ�ϰ���������
���EOAT wi?th tot�=� O�a�s߅ߗߩ߻��������oͿ�O)� S���'ϔy����� ������(�:�L�^��.Ϡѯ������ ��������*<N`˿1z ?��u�3�2C�� 2 DVhz���Ǡ�no(���/ /'/9/K/]/o/�/�/��/�v4��/�/ns&���	Advanced�/P?b?t?�?�?��?�?�?�?�?OǠ0xw�.O@OROdOvO �O�O�O�O�O�O�O_����/�/%_O_mt%�?�Mass/Center�Q
_�_ �_�_�_�_�_o!o3o�EoWoơ-32.3u��o�o�o�o�o�o �o'9K]tڶ�鿛�o_�^ ��^���1�C�U�@g�y�����\onb2to ُ����!�3�E�W��i�{�������p�w #�͏�z,��%G"0c�R�xX��R� d�v���������Я�<��c�1.5ȏ+� =�O�a�s����������Ϳ߿�� �?�@�C���)��RY� �ϸ������� ��$��6�H��-.1999W߂ߔߦ߸����� �� ��$�6�H���SžLៗ�Y�k�}��RZZ�����0�B� T�f�x�������qo�� ����,>Pb t���i�����x.����p�p�|@� Oas����� �����'/9/K/]/ o/�/�/�/�/�/�/�/ �/�(��D?*rt�ϣ?�?�?�?�? �?O!O3OEO\�n�{O �O�O�O�O�O�O�O_ _/_A_S_?|�6?�_Z?l?~?rt���_	o o-o?oQocouo�o�o ��Ə�o�o�o) ;M_q���f_�ԟ�_����\TCPVerify/&�?Method�J� \�n���������ȏڏ�쏫lDirect Entry�� ,�>�P�b�t������� ��Ο���x����=��z'��fy >������ί�����(�:�L���298.4992O�|��� ����Ŀֿ������0�Bϭ�M�C�?�/���S�e�#��?�� ���"�4�F�X�j�|���ߠ߻�	-169.1565������ ����+�=�O�a�s�����V�h�&2�)(����Ϲ�#��_@� R�d�v�����������������a951.8884��$6HZ l~������x�����Dm����9���#�W��� ����//%/7/�I/�`179.868��w/�/�/�/�/�/ �/�/??+?=?�x�3�V+�?Oa#�PN?�?�?OO1O�COUOgOyO�O�O �-.2586�O �O�O�O __$_6_H_�Z_l_~_�_O?a?�5��h?�_�?�?#�R�_=oOoaoso�o�o��o�o�o�o�o`�-2?9.4700�o  2DVhz��������_�_�S��#�_5��Z*oo?fyMean��� ����ʏ܏� ��$�6��o*[�G�t����� ����Ο�����(��:���i�'����Z)Y�k�}�axJ���� ��/�A�S�e�w��� H�Z���ѿ����� +�=�O�a�sυϗ�V����z����["����I�ntroductio��3�E�W�i�{� �ߟ߱������ߪE�� ��(�:�L�^�p�����������������9��R�t�utojog��Overview�� �������������� &8��\n�� ������" 4F��a���]��SelectT1ModeH�� / /$/6/H/Z/l/~/�/ O�/�/�/�/�/? ? 2?D?V?h?z?�?K]�o�?�?`(���E�nableTea�chPendant�?6OHOZOlO~O�O �O�O�O�O�O�/_ _ 2_D_V_h_z_�_�_�_ �_�_�_�?�?�?+oI�y$�?�Joinl`g�_�o�o�o�o�o�o �o(:�O^p ������� � �$�6��_oo{�����'Qog�ride_moՏ�����/� A�S�e�w���H���� џ�����+�=�O� a�s�����V�h���ܯ���`�HoldDe�admanSwitch��1�C�U�g� y���������ӿ忤� 	��-�?�Q�c�uχ� �ϫϽ����Ϡ�ίį�&��= ���ResetAlarm�� ~ߐߢߴ��������� � �2��V�h�z�� �����������
��.�@����[����q!M߻ą_J1@� ������	-?Q cu�F���� �);M_q ���T�f���Lo��J2-J6�*/</ N/`/r/�/�/�/�/�/ �/�??&?8?J?\? n?�?�?�?�?�?�?�0��O1O�#�cgCarȏyO�O�O�O �O�O�O�O	__-_�/ Q_c_u_�_�_�_�_�_ �_�_oo)o;o�?OVo�o�&IO��eO�o �o�o'9K] o�@_����� ��#�5�G�Y�k�}�@��No`o��ԏ��o[A�d_X��!�3�E� W�i�{�������ß՟ �����/�A�S�e� w���������ѯ㯢�ഏ��(�����_Y-Z�w���������ѿ �����+��O�a� sυϗϩϻ������� ��'����
�T�~�����_Rotation�������� �'�9�K�]�o��@� ������������#� 5�G�Y�k�}�<�N�`�0�����o��onc�! 3EWi{��� �����/A Sew��������������(/�� ���[ALastScreen�r/�/�/ �/�/�/�/�/??&? �J?\?n?�?�?�?�? �?�?�?�?O"O���/OOyO;+file/backup�d?device4O�O �O�O�O_ _2_D_V_�h_z_96Fron�t Panel �USB (UD1)�_�_�_�_�_oo�)o;oMo_oqo�o  EB�CAOaO�o���%�O�Firectories�o1 CUgy������>1�P:\\B�KUP_12-D�EC-18_01�-48-30\\ ��-�?�Q�c�u��� ������Ϗ�mJO�o�op$�B��oE�defڏ o���������ɟ۟�����#�:5Image B�B+�\�n� ��������ȯگ���X�"��m�=@'��	�k���A%gri�pperP$ToolNum.���ѿ� ����+�=�O�a�s� 6?�ϩϻ�������� �'�9�K�]�o߁�DO�R�d�������S!G��Typ�O�%�7� I�[�m����������Single �ѝ�����*�<� N�`�r������������lg�o��!�g���Comment/cmt��o��� �����#����L^p��� ���� //$/����#g/-�?���Summary*/ �/�/�/�/??+?=? O?a?s?�ϗ?�?�?�? �?�?OO'O9OKO]O�oO��@/R/�O�O�!"��/�eprogres_%_7_I_[_m_ _�_�_�_�_�?�_�_ o!o3oEoWoio{o�o�o�o�o�m�O�O�oD�",�O�M�F6�o r����������\-#�I�[� m��������Ǐُ� ���!�8/�of�(:Lss7&�Ɵ؟ ���� �2�D�V�h�'�0w�������ӯ� ��	��-�?�Q�c�u��4�F�X���|�����ss8z��,�>�P�b��tφϘϪϼ��\I�nitializ�� B�"����'� 9�K�]�o߁ߓߥ߷�@�߈������,	9>KIO/s1��a� s����������� ��,�O�D�V�h�z� ��������������
�B
���A��]�1�C�2"��� ��!3EWi (�������� //(/:/L/^/p//"A
O�/�N!��Commentv/ ??/?A?S?e?w?�? �?�?�?�_�?�?OO +O=OOOaOsO�O�O�O�O�M�/���O_�/� �OS_e_w_�_ �_�_�_�_�_�_oo �?=oOoaoso�o�o�o��o�o�o�o#g �O�O;e.o�� ������!�3� E�W�i�(o������Ï Տ�����/�A�S�e�v�JpkE���� {�����(�:�L� ^�p���������w�ܯ � ��$�6�H�Z�l� ~�������s������� �͟2�D�V�h�zό� �ϰ���������
�ɯ .�@�R�d�v߈ߚ߬� ����������׿� ��]�τ������ ������&�8�J�\� ߀������������� ��"4FXj)�;�M��(-_�!MacroNumA_  $6HZl~ ���s����/  /2/D/V/h/z/�/�/��/�/�O��/?�!���easurement�/W?i?{? �?�?�?�?�?�?�?O �/OAOSOeOwO�O�O �O�O�O�O�O_�/�/��/4_^_� %?71Weight��_�_ �_�_�_ oo$o6oHo ZoO~o�o�o�o�o�o �o�o 2DVh '_9_K_��y_�W �_���0�B�T�f� x�������moҏ��� ��,�>�P�b�t��� ������{���s� (�:�L�^�p������� ��ʯܯ� ���$�6� H�Z�l�~�������ƿ ؿ����}ߟ�S� �zόϞϰ������� ��
��.�@�R��c� �ߚ߬߾�������� �*�<�N�`�ρ�C� ��g���������&� 8�J�\�n��������� ��������"4F Xj|���q�� �����0BTf x������� /��,/>/P/b/t/�/ �/�/�/�/�/�/?� %?�I??�?�?�? �?�?�?�? OO$O6O HOZO/~O�O�O�O�O �O�O�O_ _2_D_V_ ?w_9?�_�_qO�_�_ �_
oo.o@oRodovo �o�o�okO�o�o�o *<N`r�� �g_�_�_���_&� 8�J�\�n��������� ȏڏ����o"�4�F� X�j�|�������ğ֟ ������'�Q�� x���������ү��� ��,�>�P��t��� ������ο���� (�:�L���/�A��� e������� ��$�6� H�Z�l�~ߐߢ�a��� ������� �2�D�V� h�z����oρϓ� ����.�@�R�d�v� ���������������� *<N`r�� ��������� ��G	�n���� ����/"/4/F/ W/|/�/�/�/�/�/ �/�/??0?B?T? u?7�?[�?�?�?�? OO,O>OPObOtO�O �O�O�?�O�O�O__ (_:_L_^_p_�_�_�_ e?�_�?�_�?o$o6o HoZolo~o�o�o�o�o �o�o�o�O 2DV hz������ ��_��_=��_�v� ��������Џ��� �*�<�N�r����� ����̟ޟ���&��8�J�	�k�-�������/wizard�/gripper�/steps/S?ummaryU�� ����/�A�S�e�w� ����Z���ѿ���� �+�=�O�a�sυϗ���  _��������W���ˡTCPVerifկ<�N�`� r߄ߖߨߺ������� ���&�8�J�\�n�� ������������ϐ���C�]�"�ˡG IO&ߎ������� ������0B� fx��������,>PW  �%�o�_���� �//,/>/P/b/t/ �/�/W�/�/�/�/? ?(?:?L?^?p?�?�?W�i�w��?�O "O4OFOXOjO|O�O�O �O�O�O�O�/__0_ B_T_f_x_�_�_�_�_ �_�_�_�?�?�?;o�? boto�o�o�o�o�o�o �o(:�OKp ������� � �$�6�H�oi�+o�� Oo��Ə؏���� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v�����Y���}� ߯����*�<�N�`� r���������̿޿� ���&�8�J�\�nπ� �Ϥ϶������ϫ�� ϯ1����j�|ߎߠ� ������������0� B��f�x������ ��������,�>��� _�!߃���Y������ ��(:L^p ��S����  $6HZl~� O���s�����/ / 2/D/V/h/z/�/�/�/ �/�/�/�
??.?@? R?d?v?�?�?�?�?�? �?���O9O�`O rO�O�O�O�O�O�O�O __&_8_�/\_n_�_ �_�_�_�_�_�_�_o "o4o�?OO)O�oIC��$FMR2_G�RP 1i�e�� �C�4  B�KP	 �KP�o�l�`E�ˀ �o�G[�`OH�cEP]��O���#M��-qKA��}?pIEl��`:6:N=�uq9-�}u}�A�  ��{BH��cC`}dC��=N�qB�{�uEl��d���`@UUT�UT}�R��a�>FD�>�d��>D�=��=��1U�op�H�$:��=:���:.�	:sf�:�Uf1���}� ����ۏ���8�KW�b_CFG j�kT C��������J�NO �j�F236039� 9737K�RM�_CHKTYP  �aKP�`�`�`�a�ROM��_MIN\��KS��+���p]X�`SSBZ�k�e �f�X�KUO�x���P�TP�_DEF_OW � KT�c��IR�COM�����$G�ENOVRD_D�O �VQݭTHR� � d��d�_E�NBϯ �RA�VC�clA�L�� ��f��`�}�EӤ�G
��F�/lG�,��t���KR�`�!��v���r���C�OU�`r�l� KP�h���e<�(�[5�ۿ-�^������������]�^���<,!�������n"����C���'c�>Dj�pKQC�B���W������B�`��B��a���i ɑ�.D�SMT�csQ��`�N����$HAPT�IC_CNT 2�t�e[�
!��o�@W�KSs<xҷA�KS��x�C��s2x�I��KS���H�m��s^@x�E��ۖ���ȹKS�6&x�G���KPZ�pz�7q��KS!�Z�FEAT  g�Z�� <�8��B�8T�c�X�OST_�\�s1u�iM��V_k 	������2KV��HYe��� $�6�H�HZ �y�����������f�	ano?nymous��(:L ���� �����h��� Z�7I[m��� ������/Vh z��{/��/�/�/ �/�/.??/?A?S? v/���?�?�?�?�? */</N/+Ob?OO�/sO �O�O�O�/�O�O�O_ _8O9_�?]_o_�_�_ �_�?�?O"O$_�_XO 5oGoYoko}o�O�o�o �o�o�ooB_T_1C Ugy�_�_�_��o �,o	��-�?�Q�� u��������Ϗ� ��)�;����� ��̏�˟ݟ��� Z�7�I�[�m����؏ �ǯٯ����V�h� z�����{�����ÿ տ�.���/�A�d� RϬ��ϛϭϿ�����w�Eb�1v���  P!e�#�����N�=�r�5ߖ�Y� ��}��ߡ������8� ��\���C��g�y� �������"���F�	� �|�?���c������� ����Bf) �M�q��� �,�Pt7I��m����Q�UICC0��!�11.200.�@!&/)1O/+/!  @/R/!2�/{/���/!ROUTER�/�/!
?$� ?~�PCJOG??�?!192.�168510�/#C�AMPRT�?k?!�51�0�?�6RT�?�?�?-O��NAM�E ! �!R�OBO�?5OS_C�FG 1u � ��Aut�o-starte�d6�FTPA� �AX�Z��O��_'_9_ K_]_���_�_�_�_�O �_n_�_o#o5oGo� �O�O�O�o�_�O�o�o �o�_BTfx ��o/����� ��1�C�U�����o ����Ώ����(� :�L�^���������� ʟܟ�5�G�Y�6�m� Z���~�������{�د ���� �C�ů?�h� z���������	��-� /��c�@�R�d�vψ� O��Ͼ�������ϙ� *�<�N�`�r߄�˿ݿ ������7��&�8� J��������� ��m����"�4�F��� �߱������������ ����BTfx ���/���� a�s���3���� ������/(/ :/L/op//�/�/�/��/�/pOD@_ERR� wNJ�/�&PDUSIZ  | �^��4>,5W�RD ?�E^��  guest|&l?~?�?�?��?�?=DSCDMN�GRP 2x�E;0�^| �wd|&KD	P01.00 8C�   A  �%  

@��?@}D�9 �������������hg@1g@�����XSM  �~?G�  �P��SO�ygG�E���R���{O+�?@�@�D�0k
�D�O�{g@U��@-w@�k@ew@���O�+X�I0�+Sy*d7OIO[OmO�;__GROU�0y9@�2	�1.C�XQUPD  Z�5�T�PTY�`�=� TTP_A�UTH 1z;� <!iPen'dan�7Hn�/VP� !KAREGL:*HoQo|'nb�KCxo�o^op`�VISION SET�P�o�o�g�o 'mcK9c]�������~dCTRL {=&BD|!�x $�F�FF9E3�\�FRS:DEFA�ULTV�FA�NUC Web �Servery*
 ZdT?f4�|̏ޏ�����&��$WR_C�ONFIG |��; oV��!ID�L_CPU_PC�u�|!B�_�� �A)���MIN|��D1 ?3倐?GNR_IO1:2�| 8��NPT_S_IM_DOΖ6��STAL_S�CRNΖ ��XI�NTPMODNT�OL�؛��RTY��ݖ�``ENB���R|�OLNK 1};h0�����į֯������MA�STE͐�^��SL?AVE ~?;��RAMCACHE�*�"�OaO_CF1Gl�����UO`n�~��CMT_OPu�8В:³YCLk����o�_ASG 1�7F1
 �1�C� U�g�yϋϝϯ����������	����NU�M939
��IP�i�{�RTRY_C�NͿ����Q93���b5 �������J��\0��\0��P_ME�MBERS 2���97P $�������}��(逐RC�A_ACC 2���[  QfN�� j{ �� &� 6�u��15Bo`v�"�� ~� 8�| �2�� �3��X�B�UF001 2���[= ��u3�V����u4�u4  ��u5�u5��� u�1u�� �@u�3uP��`u:u]:|!tBtp�  �� @	� `u9u�9�u7u7| ��u8u4A�u6u�6| �� u2mu�� 	�@y��`Y��q��y��u18�<Hp��	`k�x�C��1h �Hh��(�F!/`�u10�DA��u2�_A��u3T� X��u=u=7P� :i���@u o`�`a��	�`c��):��� � u3��u1;�{�u2p�3��C �C91NUNYnY�Y�Y��,)  ,)�� y�@u1a'\н��3����0�8��u�Pu+0�H�P�� �����2�������ns����#�5�G��Y�k�}�����XQ���@�4���X�����7 >���d(��?`{5���r�p��`<����cП@���Gn�/0HD�7I[m� y\�������3��(2 2!HQ(-2a"6 -2AHSLOHRYHR a�loHRyHRQ" �d��d��d��d� �"��d���d��4���2 :4���2
4���2���2 ��2*4!�b�4!�b ! �b HQ0!5B4/ �@I"�@�4X#_@:4h#  p#w@y"w@�"w@ �"w@�"� � �B��  
4�#� JD�#� �"�24��DX䊱2���]14�<�HQHP<�HP+T.QВX�HIuS�↲[ �v�� 2020-1'1-0�3{����_��_�_�A !  �|3�_�_�_
oo.nQ�g9hXt3yT9? %  ?.ouo �o�o�o�o�o�o�o�<bf�`h_zS��-�1PJ��-  M}�� # * {�R6P(Qt� ��|0' : QtHQt���,RXQt`QthQtp�QtxQt�Qt�Qt��Qt�Qt�Qt�Qt��Qt���4 �`� )  EQe�zd3y_x�Pp .� Xr;^r7�|0��P  / >xp!  7������~ , ��p+�.Q=�Dd08-2�1�:Hp_p��� !�3�E�W�i�{������P�4�؅5-2�\31w6Qd��ϒHp;��bPpϒXp0.�Q�B6P4�
��!�3�E�W�i����v���B�0x:�`Ԙ6`@[�Pp��ZXp��a� � 9 |26P � " +xp9 ^ ��ߒd�ߒl�ϒt�ˢ(|�ˢ��8F�]���D���`��ˢ��P�	���_��ˢ�p�	^�p;qK�pߒCY� �R_d_揬���п�Z&  >ۿ��*�<�N�<oNn*�p�Њ� �Ϯ����������ߨ,�,|1.�P��2� 
 SHp0:�O�Pr= Xrz�� / ' $|0;�� <��xp��\���d���  ��t���|��҄��� ���Ҕ��Ҝ��Ҥ���଀�Ҵ����p, S G�p��E�p.\�X���� �#4���� 7 	|0�Wp# 'k�Axp-ƀI�߷���������(���pp�N�p+�rՏp0����� R 7�I�[�m�������� ����Ǘ�Ԓ�Hp�Ҡ��Xp��� #�P9
��(``A��:L^�p������6r��a����Pp9�Xp��� ��|0�ҕ�;,��͠ ��͠���|������ � \��͠��5� �������p�W�  �p CY� w��������Yt /'/9/`K/]/o/]�o�9/ �/�/�/�/??%?7?�I?7߶��c Q� n1s�3 �4(^�40 q Q8�4U@�4H�4P�4X�4U`�4h�4p�4x�4U��4��4��4��4ՠ�4��4��4� r Q�`�#��A�W�4yB�0yB�0^�4�2�0�2�0�2�0 �2�0�2�0�2�0�2�0 �2�0�2@�2
@�2@ �2@�2"@�2*@�22@��2:@�2��TO-wxC�xCY_k_}_�_�_�_ �_�_����z8U�4b �0b�0b�0V�49b4�T_Yoko}o�o�oP�o��z8,�4-�4/�44�0�"�0�"�0�"�0�"�0:�4ϑ�1 ���0���0���0pr�0D���0F�4��BJDT}r@MDO&DQ.D�S6Dbh�I_CF�G 2�� H�
Cycle �Time!B�usy'Id9l�r�tmi�2'=�Up�v�q�Read�w�Dow������sCoun�!	ONum �r�s�|+䂍 Z�h�PROmG�r�����)/softp�art/genl�ink?curr�ent=menu�page,1133,������/�
��"h�SDT_IS�OLC  ����;��$J23�_DSP_ENB�  e����IN�C ���#s�A�u�? �=���<�#�
r�͙:�oi�u� �$�+��OB��C��������E�G_GROUP� 1�e��< ���͑~)��
3�?(��Я�!� ��/��S�e�w����'�=�G_IN_AUT�pT������POSREM�_�K�ANJI_MAS�K�׺KAREL?MON ����"yN�g�yϋϝϯ�(��%²������$���쿢�KCL_�LǰNU�p�$�KEYLOGGING�0���������LANGUAGE� �m���DEFAULT� {ѰqLD�q�@�����F�����G��َ�����3 ��� � '�g  �[���>�L��;��
$�(U�T1:\��D�  F�S�e�w�������������(
FRA:\RSCH2����LN_DISP �����㯹ԟOCTOL��!D�z��n�ɑ��GBO_OK ���d��������	 -?Qcs����	a	���ٍ�H���<�Ñ��_BUF�F 2�e� �2���M�0 �L^����� ��� /-/$/6/H/�Z/�/~/�/�/���DCS ���ё[0�	��sW����C+��x�]�6Bཔ|��%?�  A��>���A���>
����� IO 2��� �p�?�p���?�?�?�?�?�?�? O$O4OFOXOlO|O�O �O�O�O�O�O�O__�0_D_���ER_ITMb�d���_�_ �_�_�_�_	oo-o?o Qocouo�o�o�o�o�o��o�ok9tPSEVtΰ��nVTYPb���_m�}�R�ST$��%SCRN�_FL 2�}=������)�;�M�_�q��TP:�b�\r}��NGNAM�����m��$UPS`�G�I�p�����_�LOADJ�G �%��%J%qTU�P	�RA#�/���MAXUALRM!�,б� 瞕
E��'_PR�а ��E�Cc����k7x��k�P 2���� �$	���
ΰ�ΰ#������$� �!�Z��H���t��� �����ί��+�=�  �a�L���h�z����� ߿ʿ����9�$�]� @�Rϓ�~ϷϢ����� �����5��*�k�V� ��z߳��ߨ������ ���C�.�g�R��� ������������� ?�*�c�u�X������� ��������;M�0q\�>�DBG?DEF ���������� _LDXD�ISAˀ���1E�E�MO_APŀE {?��
 � ��0BTfx���E�FRQ_CF�G ����AM ��@����<���d%�/��ؒ���*T /V" **: _"��R/d(����/�/ �/�/�/�/�/?5?� ��^?TPO?�?s<�=�<,(3?�?���?O�? +OO<OaOHO�OlO�O �O�O�O�O__�O9_~;�ISC 1���E  ��?�_���_���_�_�_E_WR_M?STR �-}e�SCD 1�� �_fo�_�ouo�o�o�o �o�o�o,P; t_������ ���:�%�7�p�[� �������܏Ǐ�� ��6�!�Z�E�~�i��� ����؟ß��� �� D�/�T�z�e�����¯ ���ѯ
����@�+� d�O���s�������� Ϳ��*��N�9�r�6oMK��&m����$MLTARM���9'�� �x3� ���į ME�TPU� R���.iNDSP_AD�COL�� �CM�NT1� $�FN�M�Q�"�FSTLI8r�c�` �&n����������$�POS�CF��\�PRP�MP���ST/�1��&k 4�#�
 a�v1a�q��]��� ������������A� #�5�w�Y�k������������$�SING_�CHK  u�$oMODA��_[��˯�DEV }	�
	MC:Q�HSIZE�P��TASK %��
%$123456789 ��TRIG 1�&k l��~9M~=�YP�~53�EM_INF� 1�9+`)�AT&FV0E�0R�)�E0�V1&A3&B1�&D2&S0&C�1S0=�)A#TZ�/$H!/I/�=q/ (Ay/�/\/�/�/�/�/ � ?� ��	/z?-/�?�/�? �?�/�?�?O.OORO ??�O;?M?_?�O�? �?_=O*_�O�?`__ �_k_�_�_mO�_�O�O �O�O8o�O\o�_mo�o E_�oqo�o�o�o�_ �_F�_oo��So ��o���o��B� )�f�x�+��Oas �����,�c�P���t�/�������ΟJN�ITOR��G ?�e   	EOXEC1i��2�3�4�5�� �U7�8�9i�� ��|��|�"�|�.�|� :�|�F�|�R�|�^�|�Pj�|�v�|�2��2��U2��2��2��2��U2˨2ר2�2凞3��3��3"�R�_GRP_SV �1�� (m����	���jv��
�e��&|��x�����Lƨ_Dm��׳IO/N_DB' �+c�_  �c��@Z��%��c�h@ĐN ��J%�)����-ud1: RSCH\ݟ�ϰ�"��PL_NAME �!����!�R-2000iC�/125L, H�andlingT�ool  \�#�R�R2�� 1�?�(�@��R� d��'�9�K� ]�o߁ߓߥ߷����� �����#�5�G�Y�k�}���<2#����� ����&�8�J�\�n�<<����������� ��(:L^��~|�  ���  ��  ���  A�  �B� T� ���
� �� ���  ���� � B� z�� $�C��C��P� E;� E�@ D�����D�� ��� ��� 1 ��
E�):>g+E(� :9Z�H�%Z!fn/W}��Y "JJ� =��і�>>�+��f(#�P0'%��(/ 2!&!F!b%J!%2%F%�F!&!%f6)�%J!m� N+2%J!&�!��J2(��$I"�,1& S�)?$?0'� �� a2��h?n1b1F%n?�3F!�� f&!�=�g� �3�1f?�3��`�3�?�6Fp� E"B�?�3�4F�?}6>BO|7�bO��N� E$E��LE�������  � �O�K��d�C�D�O Y�O"_�0W�@��B]S��W�%n__�_KV X�X�_�ZAp� ��S�����_�_	o�W��P��TB�i����Wogl���U	`�_�o�o�o}a:��oA���o�o~ ;`\�)r�=f�_O:w |�l~{�_�X���������R�� �1���R��bl�6 Ē��� @�%?|� v���?��<v���@�6�Z1�v�)�;�	l��	�  ~�� �,^��|������ � s? � � �䂱��K�l,K����K��2KI+��KG0�K �U�����O=���@�6@ t�@?�X@I�b�������N�����
��ՙ��G��_�����v�~1a��k�ô� �"���  �X��ￒ4������r���  ������bW|��>�T���f�����	'�� � ��I� �  ��Q��:�ÈƯÈ�=���ޥ*�@����`��*�`��e4��[�p�  �'t���S���?��ab���^���C��MB� C4� ��B"tʱ����}�α*�������B�P�*u�m&p�F� ��k�	���zϳϞ�����5~ �����.�� ,0�:�d�  ��?�fafA_$�6��� w`�k�}�+�80��ߡ�?%�R�����(0���P�����΃΄8������Qa;�x5;���0;�i;��du;�t�<�!���C�R߄��`���&p?fff?��?&��Nd@���A#��@�o[��0��{��� v���t���d纄U�*� �N�9�r�]�������`������0���F.p ��,��P��q��C4�?EtPC�3�1�3̓��< '`K]���` �����g-/�T/ �x/�/�/�/M��/�/�o/?�/,??P?;?��aA�x4�P�R�?A�J?�?F8A�/C<?Ƀ��?�?OO0��m���W0OC�T��` Ca-O*�4���0�1�Ab�ܮ����bC@_;CL�n�BA��Q�>V�.È�����Y�?\���
}OOc���Q��hQ��@�G�B=�
�?h���O/`�����W���ɰ��B/
=�����Ɗ=2MK��=�J6XLI��H�Y
H}���A�12ML��jLL�PBhH:��H�K�n_�P	b�L �2J���H��H+UZBu2O�__�_ 	o�_-ooQo<ouo`o �o�o�o�o�o�o�o ;&8q\�� �������7� "�[�F��j������� ُď���!��E�0� U�{�f�����ß��� ҟ����A�,�e�P� ��t��������ί���Gϭ�� C�a�?;� Ĉ�y�]�d�CVF酿⌿�I[Կ�@��yKտؿ� 
E��� �ƿK��@(�A�_3�hM����~�����N��nπϪ�3�lC��ϬϺ¢������ϰt�.3礁}���k����q'�3�JJ ��^�L߂�pߦߔ�J�5P>�P������T��7�"�[�F�A�a�h�����{��<����  fU��� %��I�4�m����������������
���)Z,  ( 5�{0HB��~����  �2 E�G!�3Ew�L���q�5cB��0w1Q�C�l@�1  @Q�L�0� k}�b��6n��}Ӥ��0�////?�@#�8E�4y�0e��4�;
 0/�/�/�/ �/�/�/�/?#?5?G?`Y?k?}?�J�2�����V{H��$MR�_CABLE 2���� Ț��T��@P@PA?� PA�1�1�  �´ �0C�06!O4>�B����rS� ��6!�K�p(� ������?�6�,  ��� ( l6#N��/HB���)x t� BR�e�BZx,O�>L<N@` �L��D��B�%l�hB�J� .� BC�͸�] �E�?�3�O���O��O �O__ _�_�_V_�_ z_�_�_�_�_�_�_o 
oo�o|oRo�o�dE���  B���t�o�o
q��B���y�a��� ������`�� ��ՠ��@���������7p�;p�?p� ����@�����W�7p�Kp�Op���3083�/11�l�3OM ���9���K� i H��%% 23456�78901��u ����q6 �6 ;�6 6!
�w�m�not sen�t *K�6!�W���TESTF�ECSALGR ' eg�;d��a!2�
��� ��ЭD��3�l��ŏ׏� 9�UD1:\ma�intenances.xmYD,��k�p*�DEF�AULT��2GR�P 2��z  �p  ���d�6&  �%!1�st clean�ing of c�ont. vG�i�lation 56��ԓ�@ޑ��+�a��"�4�F���m��Gw� %ޮ�mech��cal checkW�/  ���C ������֯�����[�w�o���rol�ler��������ů������п�1��Basic quarterlyD�W�i��,��V�h�z��Ϟ�)�Mw���6 "8��6 �����M�"�4�F�Xߧ�6!%C;����ϸ��������
��k�}��Grease �bal�r buCsh+��}����@�������/�A�C���geu�.L�t�yN��  3d�2� :�A��	��n�����(����}�
�gG��6&f���-6 ���]�2DVhzz}�
�cabl��6"���@���
!�,>� ������������/}�Ov�erhau�ϕ�@B  x�J!Q/���~/�/�/�/�/�A$o/�/�h�o? m/ B?T?f?x?�?�/�?�/ ?!?�?OO,O>OPO �?tO�?�?�?�O�O�O �O_SO�O:_�O)_�O �_�_�_�_�__�_ o O_$os_HoZolo~o�o �_�ooo�o9o  2DV�oz�o�o� �o���
��k@� ��v��������Џ �1��U�g�<���`� r���������̟�-� �Q�&�8�J�\�n��� ����������� "�4���X�����˯�� ��Ŀֿ�7����m� ϑ�f�xϊϜϮ��� ����3��W�,�>�P� b�t��Ϙ�������� ����(�:��^�� �ߔ��߸������� � O�$�s��Z���~��� ���������9�K�  o�DVhz���� ���5
.@ R�v��������//�\	 T/I/[/m/��/� �+�-�/�/�/�/�/�/ <???V?H?�?x?j? |?�?�?�?�?�?8OO ORODO�OtOfOxO�Op�O�O�O\ ̼�?�  @\ z/Q_c_u_\=_�_��_�_\*�_** QV�P�Oo,o�>o oboto�o�o�����_�o�o�o �o1CU�o�o�o) ����	��-� w��u������m� Ϗ��=�O�a���M� _�q�3����������\\�$MR_HIST 2�U}�� 
 \d�$ 2345678901$�,���R#�9]����L�~� [ݯ����ʯ7�I� [��$�r�����l�ٿ �����ƿ3��W�i�  ύ�Dϱ���z��Ϟ� ����A���e�w�.����Q� �SKCFM�AP  U���R��Q���߳�ONREL  ��������EXCFENB��q
�Ӳ��FNC���JOGOVLI�M��d�g��KE�Y��j�s�_P�AN�؅���RU�NZ���SFSP�DTYP>�	��S�IGN���T1M�OT\����_C�E_GRP 1�U���4 �_h� Q�U���������x��� ������?��4u ,��b��� �)�"_�� |�p���/����PD_THRS�HD  Q�F�@ )�QZ_ED�IT������TCO�M_CFG 1����!�/�/�/ 
�p!_ARC_����I�T_MN_M�ODE���)�U?AP_CPL�/-��NOCHECK {?�� �� M?_?q?�?�?�?�? �?�?�?OO%O7OIO�[O��NO_WAI�T_L��e'/�OD�RDSP�#��)�O�FFSET_CAqR[ �/�FDIS�O��CS_A� ARK���f)OPEN_FILE�@��!f&� �OPTION_I�O{��QPM_PRoG %��%$�_l�_-SWOP�?�;��  ���U�����  �Ј ��Q��P'�Q	 чQ��QQ�zD���@RG_DSBL'  ����No���ORIENTT�O��?"C�����A� �BUT_SIMK_DYW�����@�V�@LCT �T����Q��$dQ��Z�dQ��b�c_PEqX� �O�dRAT�'� d)��d�@UP� ��m�!ݐ��QcI��y�$P�ARAM28��(�@�c�`/��� �%�7�I�[�m���� ����Ǐُ����!�3�E�Q�2�t����� ����Ο�����Q�<c�@�R�d�v����� ����Я�����������O��  ���  ��  A��  BC�[ B��{s3�H7���  ��?�>�BJC�zC��z`yaQ��P E;� ENE D����M�Dn������n������  ������E���Ѳ�gӳE(�ȳ��Z��Z�Ͷ�ɲ��/��%�2�B��ʱ���b�Ȳ�>̅Ζh{��汜Ӱ����3�P���ū����� ����
�����������@�������2���m��NӰ����ε^т��@�ȕ������� Bٮ�̳���ǂ�}���	�����
����<���������:�چ�� l�n��l���`��~�h�Fp �Eʰ����v�F 3�%����$炱
�4�+�0�&B�g�y��d#����������J�J�-W%P�@���`4^T
Apz?��g����q�[�� ��B�Z��2 �P�mB3	`HBTf%:�o�a����3 B�`�Z�� 2��Ia/&+(I/  /m//j/�/�/�/�F��r�pO7p1�!��(!���t>0l6!dA`_�� @��?>�>"1��?m@"1�xb�˴�"�P>;��	l22	�P *0� �,^L0�M0k0�� �� s � � ���2� H��9H��H��H`��H^yH�R�,hW��?�<� �C�PB�C�ʰC40D;0O�#�9W�� _��k��}`�ʰ�>A"O4OFO�#�B<ߟ��KA��)O�"j��OK@����C�'$/�?��? Q��V�/0_�%	'�� � NRI� �  ��MJ=���r_�[R@�_�P�N"a�_D8["b/�O�'N�`o  '�`4d�1[@B:�B}`
BoOAoSo} -�  }�
A*�8��`�>�B�&B� �f����Q�e ���/�/;&_J\pOU50`P�u�a.�u ,KB:z�L2��1�D�?�ff0����t ��)�[q8K@?�M�?���.1Rz(K@{�P ���y�1z3z4�Sj�����Zq;�x5;���0;�i;��du;�t�<!C�ڲ?��04�S|22�?fff?�P�?&,�Wt@���A#B�@�o[J�KI�b'���[p"5 �� 7���f4�֟�� ����	�B�-�f�x� c�������ү����m�������P��E C	�۴rᲂ?����� Ŀ���ӿ���	�B� -�f�/�ϕ�W�M?� ��7� �s�$�6�H�Z� ��o߁�ߴߟ�����4�����A�$� �6�C��[���텹���?�؉����l��KI�رS�W���C� p�` Ca����ʣ俣��F�@�I�Zn��bC�@_;CLn�B�A�Q�>�V��È�����Y�\���
)�����Q���hQ�@�G��B=�
?h��â�� ��W����ɰ�B/�
=�������=JMK�=�J�6XLI�H��Y
H}��A��1JML�j�LLPBh�H:��HK��, 	bL ��2J��H���H+UZBu����|��� ���!1WB {f������ �//A/,/e/P/�/ t/�/�/�/�/�/?�/ +??O?:?L?�?p?�? �?�?�?�?�?O'OO KO6OoOZO�O~O�O�O �O�O�O_�O5_ _Y_�D_i_�_z_�_�YG�y��_�_ C�a3�>�_ Ĉ��	ooOCVF�1o8o���<�o�P��K�o�o� 
E�o�oro�oz�P(�Q�_�h�o沁��*u�U�N���,��3lC�8FXfr��r���t�.3��}���|k���q'�3�JJ�}�y
�@�.��R�@�{�P�	P�����ϭ� ��0�Ώ������M�8�`�{]�l��q  fU��H�џ���� �������L�:�p�^���v�������ƫ)�ZƯد  ( 5�'����<�*�`��N�����  2 �E�����E�L�n����q��B�0�,#��PC��0��@�_��
��.�@�R�'�����ϟϱ���L�ϧ�?��ç���%���}�v��
 ��?�Q�c�u߇� �߽߫����������)��y���n{V{�H��$PARA�M_MENU ?��u� � DEF�PULS�l	W�AITTMOUTލ�RCV�� �SHELL_W�RK.$CUR_oSTYL�`���OPT���PTB�����C��R_DECSN��u� �B�T� f������������������,>gb�S�SREL_ID � �u���vUS�E_PROG �%q�%c�wCC�R�����y��_H�OST !q�!��
T���9� ;u�_TGIME���b�?GDEBUG� q��wGINP_FLcMS�`��TR���PGA� ��|�+CH��TY+PEn�z�b\ �/�/�/�/�/?�/? "?K?F?X?j?�?�?�? �?�?�?�?�?#OO0O BOkOfOxO�O�O�O�O��O�O�O__C_�W�ORD ?	q�
? 	PR��c�MAI?��bSU�~STE\�c?Xs	��RCOL�eh�Y�_@&L�  �p՜�`��d�TR�ACECTL 1��u{� �|�o p�� � ��|���:d	f_DT Q��u_`�$`D � Wu ��l`�pd�pac���b7a�a Ђb0 �bЂb	�rbT��rb�pd�pd�pdU�pd�pd�pd�pdU�pd�pd�pd�pbE�cp�bp�bp�bpp�bp�cE tUpd�pd�pd�pdT��rb�pd�pd�pdU�pd�pd�pd�pdu�pd�pb\ !pb_ �t�t߰�rU�t�tpb^tW^ �t�t�t)�t�u�t�t-�T�rs_t_&t@t�@t@N�/s@6t@��d@*�Q��s@�@+ P�P�P�� RR�P��@�@�tU@�t@�t@�t@�tU@�t@&�@.�@6�W@ P�P�P��ӰR��s@ "P�#�P�$P�%P�&P�'�P�(P�)P�1P�2�P���R�4P�5P�6�P���R�UP�VP�s�P�tP�u�g��tg�tg&�g.�g�6�g�g&�gn�g�v�g~�g *�+�蔟�g��g��g 7�8�����@&�ꒅ ꒋ��F�T��H�I�J�PQ ��P�M�g�Uh�i�j�k�Ul�m�n�o蔑p�Ű꒗�t/�\�6�u>�utu&tuJ.tu6tu�fGsuNv�	pd��u�tu�u���u��u��u��u���u�u�u�tu��tu�tu�tu�tu��tu&�u��u6�u*�u&�u.�u>��sUuF�uN�uV�u^�uuf�un�u �pdU�pd�pd�pd�pd)�pahbC&tC�c�' ��?�Ct�� ����������/�A� S�e�w߉ߛ߭߿��� ������+�=�O�a� s����������� ��'�9�K�]�o��� �������������� #5GYk}�� �����1 CUgy���� ���	//-/?/Q/ c/u/�/�/�/�(ha�% �/??*?<?N?`?r? �?�?�?�?�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� �%�/>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h� zόϞϰ��������� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���� ����������&�8��J�\��$PG�TRACELEN�  c�  �_�b��x��_UP �������������x�_CFG M�����b�������� ����� ���  �����DEFSPD �����!� �x�H_�CONFIG 9ç��� b�� k dnȇ� �!�qP�b���x�IN��TRL ������8�P�ES�]�����m��x�LID������	�	LLB� 1�]	 5��B} B4M����!�f`���� << �!?�������� �-//E/c/I/[/}/ �/�/�/�/�*y? ??K?�D?�?t?�?��?�	GRP 1��2G�  ����
b�A�P�H��@B���A} D	� Ap	@r�$I4Imm ��?�PN#´�CiORKB�@�A��O{O�O�O�O�O�B?��BC5	_B_|T^>_ <�oyQ Y_�_U_�_�_�_�_�_ q_�_4o�_DojoUo@z�c�ob�
o�ooo �o�o�o>)b M�q�������b:)b�)
V�7.10beta�1 @��{@�A&�H�1=�C� CzB��O�D1� e�C��� b��� D�nw�A@ �1B M�@�1C�1 �� �!�!C�����B��0L���%���0C9RL��	�����AK33AFf?f@s33BZ�z��!A�ffA�3�3@����^�}#E�N���b� ���O��Fq���m�������
KNOW_�M  ��SoV �]
� ��oQ�c�u�Ɵ�������ϯb�,MM�3ͮ] �M�	�������:���*��Ic�$@>�� y�u���� MR*�3��T�J���b�C�cU����O�ADBANFWD�� ST�11 1�ϧ�?�4E�OAT with� tote�B@?��  �L�3�3F���G��3F��fc��]�nof�Ms� �����Iش���� �������/�a�S� eߪ߉ߛ��߿���� ���L�c�<�2G��}4/�  �<��X��03n����<�A4��������<�5�&�8�J�<�6g�y�����<�7��������<��81C<�MA�'�-Dk��OV_LD  c3���>�PARNUM  J��\�39ǷSCH�	 �
�IW5�iUPD��dE���_CM�P_��� K�6�'�3��ER_CHK���3������RSư*��1_M�O'�J(_7/_�_R�ES_GF��c
 ���/d=�/�/�/�/? ??I?<?m?`?�?�?@�?�?��#m��,�/ �?�%���?OO�#� 3OROWO�#f�rO�O�O �#��O�O�O�# �O __�#_ /_N_S_�"�V 1�J�/���P�`M"THR_INRư��3Žd�VMASS�_ �Z�WMN�_cMO�N_QUEUE ��J�3�[ � *_�N�U!Nf:h�QcENDVat/piEcXEope�BE~`|`oQcOPTIO]g�}+T`PROGRAoM %4j%S`��_8RbTASK_�I��nOCFG ��4o�([pDA�TA���d{@�v2+���
�� �;�M�_�q�������ˏݏ�zINFO��ը}(�ȓ�0�B� T�f�x���������ҟ �����,�>�P�b��t������ �֨| ��9ZqPK_^qq�dy �ۦENB� H꭮�
�2�%�G^q�2�� X,{		!=���q�����$U�!������T֧_EDIT� �d߿�WtW�ERFL�h�S9�RGADJ �κ/A�  <�?[ H���Q �Ta��_�?�A�z���q<��)%DIAG���Ϻ�	_¸��2�j��	HK`l���RBp>���UU@x��*z,�/.� **:7�P'�9�Yߺ�P>����@�u�ߴب�Yz�8>��:�߬��߸��ߺQ�PA�����g�%�7� L�v�����t�������r����>���v����A P
�^�X�j������� ������P��L60 B�f����( �$�>� zt� /���� �l//h/R/L/^/�/ �/�/�/�/�/D?�/@? *?$?6?�?Z?�?�?�? �?O�?OO�?O�O 2O�OnOhOzO�O�O�O�O�O�O�	w�_�xo_�_�T�t$ �_��[�_�_�_o-oZ�P?REF �j����
 �IORI�TY�gն�$�MP�DSP�a����gU�TFv��ODUC-TCqκ0o��;OG��_TG�Hr�Һ�bHIBIT_�DO�{TOEN�T 1�λ (�!AF_INE��`epw!tc�Љ�{!ud���~!icmX�]��bXYc��μ;��)� D�$�6����_�B�N� ��r��������̏	� ��-�?�&�c�J�����I*�cc��j���%G_xݟ�yb>�%�"օD�/N�˟@�����������,  �``Ρ���������
e�0�Z0����#��5����ENHA?NCE 㺝��AЫd/���|��fId��Qocc�$�PO�RT_NUM�c��e$�_CA/RTRE{�	�ZSKSTA�g2{S�LGSbp�	����Ù`Unothing��zόϞ��7k>�TEMP ���i��?Ub�_a_seibano � o�C�.�g�Rߋ� v߯ߚ��߾���	��� -��Q�<�u�`��� �����������;� &�8�q�\��������� ��������7"[ Fj�����|���VERSI�`��g. di�sable����S�AVE ��j	�2670H72%2��!������ 	��bA_+/�ce,/U/g/y/�/�*D,��/˭�K_p 1�	��w ��:�
W?+?WB`URG�ET�Bp+~�qWF W0'q�dj��fW^px4��a��WRUP_DELAY ���k5R_HOT �%fV�a���?�5R_?NORMAL�8�bx�?<OGSEMIO�AO�O@aQSKIP�#���3x��O� �O�O_�M^]<_lS@_ f_x_�_P_�_�_�_�_ �_�_�_,ooPoboto :o�o�o�o�o�o�o�o :L^$6� ����� ����6�H�Z�K3RA����Kh�H��t�_PA�RAM�A2�K; @g�@`�&j�W2Cu��BÁ�C�&ձBt�BT�IFy4�RCVT�MOU&����t�DCR�#�I� ��AE����EDE܅�vD��C���OB��(��Gţ����Љ�	����9�Ú?�A�z�O���_ ;�x5;���0;�i;��du;�t�<!��ذ���&���J�\�n����������ȯگ������R�DIO_TYPE�  �-��EDV��T_x����X��BH�#E��j����nz� ��B�� ��Ϻ�������=� (�пn�mO��$_��� ���������4�"�X� Bׄω��P߲ߠ��� ������
���T�v� {�ߜ�6�������� ����>�`�e���6� ��2����������� :\�a��B� ���� �$F K]~��� ���� /BG/f (/z/h/�/�/�/�/�/��/�/,/R/C?�j�I�NT 2��9���4�G;� �?�;�x ��?-�f�0 �? �;?O�/OO/OeO SO�OoO�O�O�O�O�O _�O�O=_+_a_O_�_ �_}_�_�_�_�_oo �_9o'o]oKo�o�oyo �o�o�o�o�o�o5�#Yf�EFPOS�1 1�9� � xAT HGOME��Ճ��(�1���z��lu��
�Ż�����x�����(�=�5�}@N���=1?����?�H�3�l��ABO�VE LEFT JACKP(�Ň���+^��H�~�F�f#���4���+�ɏ���|�~���ڍ@���z���RIG�H����,^�@I����G�*;��"y��nʿ�ʏ܏� �"�\���X�џl��������+��O��E�O�pchangeO pos�w�g���?��x=�̅��<<!H����%?�N�p�����MAf0� 1��d��ɾ�I�/���E��<Lu'����������ί��2��e����>g�࿊H��<ǘ���x4���"�8�F���3c��f��ʣ���
ٿ5S��;j{�?3k����������At Palle?t Stop餡��o����>�����=�9)�D��t8>[����(�6�H�a���p����ҽվQ@����8xv�տ�T[��^���ϠϮ���ٴ��q���d��>	�
��
Ee�b����謹�����&�8� 4|�r�&��=�����6K�f����!�4�]�zߐߞ߰� 㡉s����69�Յg�����3����_a��!����'�p 6|�t���B�E=�E���	�I�������/���Fe j�����<�M�8� q����0��������� ����7��[m T�P�t�� 3W�{� :��p��/� A/�e/ /o/�/�/�/ Z/�/~/?�/+?=?�/ �/$?�? ?�?D?�?h? �?O�?'O�?KO�?oO 
O�O�O@ORO�O�O�O _�O5_�O?_k_V_�_<*U}u2 1�3_ E__�_�_!o'_Eo�_ ioofo�o:o�o^o�o �o�o�o�oeP �$�H�l�� �+��O��s�� � 2�l�͏��񏌏��� 9�ԏ6�o�
���.��� R�۟v�����ԟ5� � Y���}����<���ׯ r��������C�ޯ� �<�������\�忀� 	Ϥ��?�ڿc����� "ϫ�F�X�jϤ���� )���M���q��nߧ� B���f��ߊ����� ���m�X��,��P� ��t������3���W� ��{��(�:�t����� ������A��>w �6�Z�~� ��=(a��  �D��z/�'/ �K/��
/D/�/�/ �/d/�/�/?�/?G? �/k??�?*?�?�_�T3 1��_`?r?�? *OONOT?rOO�O1O �O�OgO�O�O_�O8_ �O�O�O1_�_}_�_Q_ �_u_�_�_�_4o�_Xo �_|oo�o;oMo_o�o �o�o�oB�of c�7�[�� ����b�M���!� ��E�Ώi�ˏ���(� ÏL��p���/�i� ʟ������6�џ 3�l����+���O�د s�����ѯ2��V�� z����9���Կo��� ��Ϸ�@�ۿ���9� �υϾ�Y���}�ߡ� �<���`��τ�ߨ� C�U�gߡ����&��� J���n�	�k��?��� c����������	� j�U���)���M���q� ����0��T��x %7q���� �>�;t��3�W��?�44 1��?���W/B/ {/��/:/�/^/�/�/ �/?�/A?�/e? ?? $?^?�?�?�?~?O�? +O�?(OaO�?�O O�O DO�OhOzO�O�O'__ K_�Oo_
_�_._�_�_ d_�_�_o�_5o�_�_ �_.o�ozo�oNo�oro �o�o�o1�oU�oy �8J\��� ��?��c��`��� 4���X��|������ ď��_�J������B� ˟f�ȟ���%���I� �m���,�f�ǯ�� 믆����3�ί0�i� ���(���L�տp��� ��ο/��S��w�� ��6Ϙ���l��ϐ�� ��=�������6ߗ߂� ��V���z��� �9� ��]��߁���@�R� d������#���G��� k��h���<���`������A��*S�YSTEM*��V�9.10170 �G9/18/20�19 A � � 4��#51�_T   l �$COMMEN�T $EN�ABLED  �$ATPERC�H�DOUT_T�YPE� �IN�DX��	   w 	�TOL��HOME� �
i6qw���\��  i7q�*<N`8qq������`SMSKr�  $MAX�jEN����i MOTE_CFGr? T $�$"�" �#IO �*I�, �!LOCAL_�OP�%�#STAR}T{'POWERr� m FLAG� �"�"r ,� �&$DSB_?SIGNAL�"�"?UP_CND�!"�S232�% �� ��DEV�ICEUS�#SP�E �!PARIT�Y*4OPBITS��"FLOWCON�TRH �!TIME� �"CU�0M�"A�UXTASK�"INTERFACi4�TATU�0����A0CHr 	{ t�OLD_o0�C_SW"FRE�EFROMSIZ� "� GET_DI�R�	$UPDTO_MAP "� Td wENB"EXP0JzC!`0FAUL@�EV!�RV_D�ATA�1
  �$d@E�1   =? VALUyA> �`FGRP_ ��"dA  2
 ��SC�"	� ��$ITP_vB� $NUM�@O�U�!�CTOT_A�X�1�CDSP�FJ�OGLI�3FIN�E_PCZ1�1ONED�Eo!�@�6K+@O_MIR�ATP� �TN5XAPI 0!RE_EXXP2D�A5 �.Q�"�APGmVBR�KH�11FNC�@I:!  �R#�R�B�P!@D�!�C1PBS�OC�F� N�UDU�MMY163�BS?V_CODE�!*3�FSPD_OVR4 |@�LDb	S�ORg N fFؕP2g�@OV�ESF�JjRUNMc!!SFxff�!SUFRA|j�TO�4LCHDL}YWRECOVd �@WS @�P�e�@�RO�3�QP_f` _  @� Su@�NVE� !OFSr�`C�@ "FWD.a��d*a�Q�QU�PTR�)1o!_VQFDO>QVMB_CM�!<pB�@BL_c S^r
dq2ncV�1 "@s@d�CFbG_wrXAMpS`Rp�0�u�b�_Mvp�2M�@�"�`T$C�A�@�pD�R�pHcBK!A0F�IO%q��!"�PPA	��5��E�-��u�"�bD?VC_DBG #w�@1A2w��b�!��1����s��3���`ATIEO� �1�0aU #�@�&CAB P" "@P�d1 �x!!�@_�0~0FSUBCPU2PSIN_0Hs�t�"@1D�ws�t�"�Q$HW_Cq �0S��$�|�wq
 @|@�_$UNIT�T��>��ATTRI3@���PCYCL#NE�CAۂBSFLTR_2_FI-#/9��"6!!LP[CHK�_�0SCT4SF_ƛ�F_��.���FS8!1�r��CHA=��po�r�2n�RSD�``2�Q;C1� _T�x�PROǀ6s�0EM _�@�ST\�S�|@�\�wp�DIAG~1ERAILAC��*�M�@LO�P!�VM4�BPS�B" #����sPRx�S$@ I�M�Cj�\0	�c�FUNC�R�1RINS_T$A ���m��1RA~��@; ��p��p �t��WAR�BP�CBLCUR���ǴA����ø��D�A�P���ǳ��LD@@�P"�)��A��.��)�TI:�IſA|@$CE_RIA�1V+2AF:�P91t�,�`z�T2�C/C���qqOI��9vDF_aLy ~bA�0LM�s�FA�`HRDYO,BQ�`RG.�H��4Q� 	���MULSE��3CI��P��$J�jJ,bAg<kFAN?_ALMLV)3H��WRNO�HARDH !F�P�2��2G�Ȅ1�A�U_�`0FAU��0Ra��2TO_SBR�%���@�ڛ�l�|u���MPINF�`��������REGF&NV@��VD� �NHtFL}��R$�Mʰ��3I��p|@lV�]�CMj�NFƑF ! �?pprk ;$-!$Y��A� �B�As � �eSEG���C�PF��AR�@�#�U2�S����rUAXE�GR�OB�JRED�FW�R�`�Q_#��SSYЖP��PE�SO�WR1I�`��{�ST0�C(�0�P `E��? ��)����@B���a��5\��pOTO�? �`ARY�C���˄�="�0FI{P�3$�LINK��GTH���8@T_���ar��6�BXYZ!B:
7-OFF�`��)��B�@b��r�a)0@sFI@ʐ��0*3�Tb��D_JZ1|Bb��"�������8�Bg0����2�C�!bUDU	r��]9*�TURJ�XPÈ4����X^��p�FL �`����R6���30�Bq 1J? K PM0D�U3S��-�I�:�I�	CORQ����A���wq-�xPO A�z!b�$3C�A�$'OVE!��M�0! ��8%��8%��7&�16'0$A6'@5$ANs��� 8!z���!/Pw ��! 0%!<'�%���%\#�ASERQ��	.�E�`Hd@:��$A�!|@�����������AX �c|B�������Y5� e9�e9)�d:��d:, �d:K d:� d:+d:1 �d6��a9��q9���9 ���9���9���9���9����9���9�1�9DEBUs�$n�z���ArAB��.ar#V�pr� 
�B �����Ewq�G�Q�G)� �G���G,�GK�G���G+�� z���sL�AB��o�|�G�RO���s��pB_ȡ�&{�ã� �КV��Q��U���VAND �.��$��!��g �q{��'h��6h�� NTZмcY`VE�LΡ�$ca�kf�S�ERVEY`�� i$����A�!�`�PO�bs�Ap��a؆b�!����$.�bTRQ��
�c.��`�gz�2�fX��?_  lX��qN�ERR�q�I�p8g`�$,qTOQ�$� AL�c4k�?v��G�e�%� ��aRE>
�  ,�a�e��`�"RA�q 2 d�r-���}s�`7 ��$, ͢l��S2G2�cOC����p  {C�OUNT��xsFZ�N_CFG�a 4x���T�p��p�CV�@�q�����^�� ��@M=��!Ҡ�Հ�#5!=�u�F!Ag��%u�y�X� u�Uq���d��9P����HEL7��� 5� B�_BAS�RSR�V��S��B���1hw�2*�3*�4�*�5*�6*�7*�8hw��ROO�op��f NL��AB�c� ��ACK�FIN�pT!�M�U����a����_PUt��OU�cP~���ivb��}�?6TPFWD_�KAR1q#� pREĥd��P�����QUE麠 ltЇ�IK��C� �h`�SEM�A���A���Aq�STYɔSO����DIՑ{�7�u��>7��_TM/�MA�NRQ� END���$KEYSWITCH�-��~��HEBEATM6`�PE��LE0r����P^�U,�F��-�S~�DO_HOMx��Opѽ�EF� PR�x9�0�|�֕Cx�Ox��p�qOV_M�<s�Y�IOCM����A���HK��# D�G�Urs��M��G�X FORC �WAR�·b��OM��  @��D���U��P��1(z�]�|�3z�4���b*�pO=�L`��r�OUNLO�t���ED��  �S޲PHDDN�a ��`BLOB  �^�SNPX_�AS� 0D�A�DDG�I�$SI=Zuq$VA�Pju�MULTIP�����A`� � $�Ь�� ���S7��QC,py�FRIF���pS]�oɰ��i�NF	�ODBU ^�8`zսӸ٥fw� ��IAN��������S��� � �#�IrTEm��SKGL1�T��^&)��J�SG�2�STMTdkc�P��o�BW �3�SHOWk���BANw�TPU �+�����{pV� _�GY�  � $PC��P�p�#U1FB\�P��SP��AԐ��P��VD��X�!�; �qA00d1� ��9���9���9���9�U57�67�77�87�97�A7�B7�n�9�mQ:���9�F7��0���C�����]����w�1���1��1��1��1���1��1��1��1���1��26�2C�2�P�2]�2j�2w�2���2��2��2��2���2��2��2��2*��2��36�3C��T�]�3j�3w�3��U3��3��3��3��U3��3��3��3��U3��46�4C�4P�U4]�4j�4w�4��U4��4��4��4��U4��4��4��4��U4��56�5C�5P�U5]�5j�5w�5��U5��5��5��5��U5��5��5��5��U5��66�6C�6P�U6]�6j�6w�6��U6��6��6��6��U6��6��6��6��U6��76�7C�7P�U7=I7JI7WI7dIU7qI7��7��7��U7��7��7��7��Y7���rVP\�U�b�"�¶P�
�`V��Ҏa# x $TORf������r�`�R�`ڀ�TQ_�pR��`Au�a8�ndSmC4��e5f_U��@a���YSLfp�`$ � #���$�������� ��ld��VALAU$�ߐ2�a�hF]a�ID_L���eHI��jIN�$FILE1_��d#�$��E��[cSA�q% h��P$pE_BLCK�`�1rL�:xD_CPUJy$�Jy�/��ot��Y1� �R &? � PW�p��l���qLAq�S�p��t�q�tRUN_FLG�u�t�q�t0��u�q�t�q�uH ��t��t��T22�_LI�`�'  ��G�_O��:�P_EDI��MC2���:�(B��ɲ�Eqk�,���TBC2#�) �(�$��p����:��FT����ãTDC"�pA��Q�ɀM�PÆLفTH�Ѐ����S��R�����ER�VE���ã������ *Xw -$H�LEN��0U�ãH��RA\���&\`W_aws1H��dM2��MOBq��S��ҐI�1b�a���TH��̛DEܕ��LACE�cCC��1bp�_MA	�ۖ���GTCV�=��T� >�]�S��ړ�ၥ�*��JΠA��M��f��J��!�ڕǡ�T�2������ٓ��JK�VK��� �����J���	�J�J�JJ�AAL�	�?��?�9��=�5��p�N1d�p�/���dL��__�����v��CF�+ `�PGROU�`M�����N��Ca���REQ�UIR�ƠEBU�x�D���$Tܐ2�*�E�붎�Д�,� \B`t�APPR���CLb
$K�NN>�CLO��N�S��c�ڕ
��L�- ���M׀�o���_MG�Ѩ�C#�%p�ȸ�����BRK��N�OLD�ƒ�RTM!O9����͢�J9���PA���������]�(��f���6.�7.�?��qD���.� ��o����� ��PATH�ױѧӱѐt��ӎ��-3a��S�CAx���?§�INFG�UC�����C�KUM�Y��vp�� ��a#�2��2�H�2�PAYLOA��J{2L�PR_ANρs�L�p}�y�m����R_F2LSHR���LO~�U���|���ACRL_:q ��� �e�g�H�`b�$H��%�FLE�XA���J��/ P+£����.���|A�G�0 :T� f�됷���i�h��r�����F1��0��@��ɟ۟���`E	� �-�?�Q�c�u����� 7T�����D f���̯ޯ���T�5X =a>����%� ��,�>�B�K�9�]��f�x�������J��1 �����ο�퀺PcATI󱥠EL� ���3��J�0�J�E��CTR �DT�N�Q6�HAND_VBbA�`��72 $�F2�����cSWA_EN�����3� $$M�����P���8���<� �5��6A�`j�ƈ�aI��A�̖`��A���A��@��cp��D*��D��P��G�p�ICST�ǼA�ɼAN��DY�p<����4&E�� I��������l�������P6�?�H�Q��Z�c�l�uԢ��41 �0���� q�U<p��QASYM��@`	����3"a������_�����	�d�8 )�;�M�_�q�Jx�)����c�i��V_VI�r3�hp��`V_UANY��`s.#��J�� %rSU%r��)t��6tZv ����)�
���u��2�:�  1���HR��w�5�2�qT�&N�DI���O�t>��p��6 > -BIaA-���'�J 5c5��M '0�� �p 7o � �1ME��� P��r7aT�pP�T�`� ��x����� S�o`}�����T�`��� $DUMM�Y1H�$PS_fG RF	 �p$ӆ���FLA��YP��킀�$GLB_T�0�u�x�\�8� H1T�8 X+��ւ�ST���SB}R��M21_V��T$SV_ER��1Ob`N�f�CL"�N�eA� O*��pGL�`;EW��9 4����W$Y"Z"W��頲�3AQ��`��]U��: �Nːޓ`$GIX0}=$�� 9x0��ʐ��; L���ab�}$FabE��NE+AR� NNF;�� �TANCN�QJO�G��� <	�?$JOINT�����r��MSET��=�  �E!�K� S��"���!��>� �E U�?��L?OCK_FO��1��pBGLVK3GL��TEST_XM�A���EMPw�^8	� �Р$U��F 2:�ʓ/�;��h�0ՠ/�9P�CE��|��P� $KAR�}M�sTPDRA��m�d�VEC��~�h�kIU/�<4�HEנOTOOL��V;RE��IS3��ò96Q�D ACH���E=��O�Ѐ�3>!���SI1�  �@$RAIL_B�OXE�s�RO�BO �?�s�HOWWAR-��Ѐ�ROLMۂEū!��V��!�8 ��O_F�� !s�HTML�5�q ��sGX�C�H��?p� �R
��O��@p� y�}����_OU��A 	d��+�97a!2�!Р_$PIP�N�����ݱV /�����CORDEDՠ�п�&8�XT��)�p� �O7� B D �OBSA%3ՠ^��MѼ��M�a`'1SYSM�ADR&1�px��TCH�0 C M,�EN�r]�Aܡ�_��Դ!���V�WVAS�D �� s����uPRE�V_RT`Q$E�DIT��VSHW�R�!:�������`Db�&!5�.!$HEADra�pO���a�KE����C�PSPDf�JMP�j�L�u֐R� �QEU�R��I
�S&2�Cl0NE��'1b7T'ICK�aM[�R���HN0�F @pWЭ�%n�_GP���^�STY���L�O"��������G� t 
��G��%�$���=:�S !$q g��$��9P�P��SQUg�<��aTERC|��R��TS�$H  �F��'��'g��(01O}�p�R IZ����ρPR3�܁̩���PUq+_DYO@���XS��K�v�AXIJ i�4�UR� �'2&���x֗1�� _����ET�P(ޢf��UI�F�WJ�YA�A�QÄ9��>0 ��rSR4Il���9��:�6 �2GII LAGLQGLaF^x �I^��R|C���C�Zolo~o�d�S}C
� J hs�cDS�n�SP!�&x%ATO@�2,����⿂ADDRESz��B
�SHIF�#^&�_2CH&0tѹI)��!�TU)�I��1 Kp�CUSSTO���V��I�AL���!�P
	��
��V��;U�M 	\�����I�<���W2C�C��):��l��W1�TXSCRE�EO�N�pe�TICNA�����4��q8��"�PO T��i� ��h�E��6X��X�4�RRO*PU��а`��1F��QUE��P# ��P���S����'RSM��NU<е��vaA�pS_ē�Fc qA�I�Gc�Cʢ]B��4 2O�0UE¬TQ�y��F GM�TmpLGqgU�O^z�BBL_�W��NU�R �I�!RO��-RLE�"8S%��"�7TRIGHASBRyD{��!CKGR���iUT=�hWeQWIDTH�+�E� �큭�� �UIx�EY� T�S��D�-��=BACK+�ۂ4�U�[�FO*��W�LAB6?([�I<�΢$UR+�`���Pa�HA T 8�qU�_N��"?b�b�R��Т��ˁ���+bO�!U�U��$��bPUMP�cRޢP��LUM�co� ERiV��?AIV�NE�T5VY�� GE b&��� C�W�LP�e�E��=!)�g\�
x]!
xTװ	y5{6{7{8�b��p� ?�k4��jױȡS��U�Q�USR��W <ğ�a�U��#�FO\� �PRI�m���{q�pTRIP	��m�UNDO�X�n��pP7�O�@8'�� �� Y:b�p.G V�Ti�+!L�!5�OS��J�R� B!���1�Z�������q����&�U�a1�[�z����C�b�!�OF�F��2�\6���O � 1Zs���-[s�GU��P���p-�(!7��QSUB�L�� �RTs��]��T�u���OR�}�RAU� ~�T����c�9_�Е�^ |���OWN$���$S#RC(@�@l�D����MPFI$�S!� ESP'���0���c�<�gɲ������A_� `ÀWO2������COṔ$� &�_���w���~�WA
�C���[�1��Z�?� ���C�1 �`�2SHADO�Wl ��͡_UNS�CA��ͣ�TڣDGyD�e�EGACq�l7��PG�2a:bNhSTE4Q:�Ox`��d�PE�bgVuW��qTRG� ��Ab ���0�MO�VE(C��ANG��D��؃������LIM_X̃��҃���� ı���CK��p� �����VFi ~��qVCC�M��c�2C^�RA�O�@�z�� 5�NFA�����E�a2�pG� APb��&�DE^�
1�.E��Ad� ��z�ADű͎�dcpC����DRI����j�V������� D�tMY_UBY�tE�q�z�)A���0<�@�?�OңP_�$�a�L1B�M4Q$��DEYƵ�EXP5C��MUb��X7���v@US��v �p_R�1���p� z��G�PACI� g�󑋴��؃�җ����C��RETb�!q�Rq���ҙ�e � 
i�Gk�P�29��`��	Ra���f�P�`A�Q�]�	v�HR6�SWH���P�� O�q��QA� ��EzpU�<�]�P�@��HK
A�g�`�ꏱ� ���0��EAN��Z�A`x��i���MRCV�AWh ��`O5�MA`�C�3	=��6�=�REFW_�F�1񵲸 ��pB���S���d���F���_������ 4�4D2Ҟ0#�C����Di �H�l0z�#��q�$GROU@v ��0�mE�w�dO�,!2e�@�0m08�P�f�#,!�R@� U�L��g6�CаUah�Д NT1��?�@�na��q�� LK�@
[�
na�q1��T�DDj tÀM}Di�AP_HUZ�쐰VSA��CMPB(@F\um]_t!AR�S!��X���VGF����k� �`M�pAP0�UF_&@v�/��uROKP�2�7դ`F��P��URE�RA&��RI��_I� g���������ȹ�҃�IEN��HT$#ȜPV�� ײ?��#{S�%W��'�����Á���-9��LO������#P9�\1uqN{SI�VIA_Z���0l �+PHDR{ �P$JOup�R�$Z_U�P԰-BZ_LOW �5y1�GaRӰ[AL P�W�B��1y1- \@��g�0�����m�� 0�PA�Q= �CACHc4P1�(EO1��DI�a���CJӱI�F�1pET<P�oF'$HOA`ܒ -@��öb"�FP�R`����aT�VP3�<]��B_SIZZ��D�Zg��H�1�G��|SM�PZg�IMG[��N0ADMYw�MRE�SmRWGPM��N�D����ASYNB{UF��VRTD�U��TQ�COLE_2�D״�U2܀C�U��[@Q���UECCU&�VEM�(EbnGVIRCMQ�U�S�b�Q&0LA+���(���<�AG�YR��X#YZ� ����Wj�h��!~dS�,`TE���I�Mea�VGb�cEGRABBn�Y7�;���>n����CKL�AS*@��AK@o�  �`T4�p@Ģ�ܔ$As��p A�v!��0b�#LuT� ����7��r#�Ist'��Kf��BG_LEVE����PK��Mf�6PGI<pNO7����(�x�HO���q � w�_� �P�v�S�0���RO��A�CCE��]�#�VR_c��M`$������pARE�PA��S�� }Dq�REM_B�d��p7rJMP  ��r<t�$SS�����7r[@zQ@s/  N2SoPJ6�Nڄa�LEX=vt�Ȣ����� �DDR��$��Ӡ�}�\��u2P2Fu�� i!?�V_�MV_PI�Su�T���z���j ��F�0�Z ������y��!���!���h�GAɕ��LOO~���JCB��~w�Cx���@֣PLANҲqB�r�F"SO���P\�MQ�)�Ń���S+К�P����!P�nB �!��PâT?��P�RKE�N�VAN9C���R_O�@v (B���ɳ�S��S��bR_A�� w 4R�!�ΰ��p�I ��@x h��ࢉ}1�W�OFF�v�F\`eDEA�j�
�P�PSKsDM8���� w ���@|'�ry < ��-��UMMYj2�D2��4q�CUS��U��z� $� TIT��$PR�+�OPLG�t3SFD�\�{p����P&t�p�MO"�|Ђ�K�J;���K�0Q_�E�}Ђ�X���0��@�X�S�~ x�0MSGPD_���1�`P��`�S40NB�2LNTK3�M�>4�p�C�0#���1Ҷ�'1o�XVR��b�X�T6���ZABC=�K��-�~�

AZIP�Y�Ђ�pLV�CLw��~�6:�ZMPCF�Ղ~���3��V�DMY_LN�ϰı��� �ԃ� $�A ��C�MCM^ C�CCA�RT_G�k�P8� �$Je�_�D �Ak�|�u� �� _�0R�Y�z��UX�a
�UXEUL��ap� �������������d��FTF�k�%�m�{�Z��� �˨w�5p?�Y�0D�` �� 8 $R�[PU2��EIGH��X�?(� ����8v�?�>� ��pf�q!��$B� �0}2�SHIF���RV2=�F�@��	$��6�C�0`�U�f�0��
Ks&�D6T�Rb �V�Q>�SsPHB�K� ,� Xz�������0F� �5 1 ����  x��I ���	 ��� � �gR�&�J �n�	/�-/�Q/ �u/�/"/4/n/�/�/ �/�/?�/;?�/8?q? ?�?0?�?T?�?�?�? �?�?7O"O[O�?OO �O>O�O�OtO�O�O!_ �OE_W_�O_>_�_�_ �_^_�_�_o�_oAo �_eo o�o$o�o�oZo lo�o�o+�oO�o sp�D�h� ��'����o�Z� ��.���R�ۏv�؏� ��5�ЏY��}���*� <�v�ן������� C�ޟ@�y����8��� \��������ޯ?�*� c�����"���F���� |�Ϡ�)�ĿM�_��� �Fϧϒ���f��ϊ� ߮��I���m�ߑ� ,ߵ���b�t߮���� 3���W���{��x��<��6 1�S� e����A�G�e� � ��$�����Z���~� ��+������$�p �D�h���' �K�o
�.@ R���/�5/� Y/�V/�/*/�/N/�/ r/�/�/�/�/�/U?@? y??�?8?�?\?�?�? �?O�??O�?cO�?O "O\O�O�O�O|O_�O )_�O&___�O�__�_ B_�_f_x_�_�_%oo Io�_moo�o,o�o�o bo�o�o�o3�o�o �o,�x�L�p ���/��S��w� ���6�H�Z������� ���=�؏a���^��� 2���V�ߟz������ ��]�H������@� ɯd�Ư����#���G� �k���*�d�ſ�� 鿄�Ϩ�1�̿.�g� ϋ�&ϯ�J��Ϲ���7 1��ϒ��� J�5�n�tϒ�-߶�Q� ���߇���4���X� ����Q�����q� �������T���x� ���7���[�m���� >��b���! ��W�{�( ���!�m�A �e���$/�H/ �l//�/+/=/O/�/ �/�/?�/2?�/V?�/ S?�?'?�?K?�?o?�? �?�?�?�?RO=OvOO �O5O�OYO�O�O�O_ �O<_�O`_�O__Y_ �_�_�_y_o�_&o�_ #o\o�_�oo�o?o�o couo�o�o"F�o j�)��_� ���0����)� ��u���I�ҏm����� �,�ǏP��t���� 3�E�W����ݟ��� :�՟^���[���/����S�ܯw� �����8 1߭�����w�b� ������Z��~��� ��=�ؿa����� �2� D�~�����ߞ�'��� K���H߁�ߥ�@��� d��߈ߚ߬���G�2� k���*��N���� �����1���U���� �N�������n����� ��Q��u� 4�Xj|� ;�_���� T�x/�%/�� �//j/�/>/�/b/ �/�/�/!?�/E?�/i? ?�?(?:?L?�?�?�? O�?/O�?SO�?PO�O $O�OHO�OlO�O�O�O �O�OO_:_s__�_2_ �_V_�_�_�_o�_9o �_]o�_
ooVo�o�o �ovo�o�o#�o Y �o}�<�`r ���
�C��g�� ��&�����\�叀�	��-��%�MASKW 10�'�q���Q�XNO  �`�~���MOTE � ��!�֑_CFG� ݝ
��P?L_RANGّ?��4���OWER �0�R�9�SM�_DRYPRG %0��%ڏ��X�TART J����UME_PRO�g�y���!�_EXE�C_ENB  z��5�GSPD͠���$�TDB�2�D�RMS�D�IA_OPTION*��
�7���NGoVERS������H�I_AIR7PUR(� ժ��\
�F�MT_Y�TE��ۛ9�OBOT_I/SOLC�������K�NAME����˿o�_ORD_NOUM ?��R���H722 � ��������Q�P�C_TIMEOU�T*� xQ�S23�2��1��C� �LTEACH PENDAN�X�����ُ�׀Mainte�nance CoKns��jߌ�"���ӄNo Use zݶ�|��������"�O�6�NPO�� �����3�CH_LfР	7�#�	��~p�!UD1:��zr�RX�VAIL��曵�5���SR + �����~��R_INTVAL����5�V��V�_DATA_GR�P 2��
�� D;�P%���!� ������>, bP�t���� ��(L:\ �p������ � //H/6/l/Z/�/ ~/�/�/�/�/�/?�/ 2? ?V?D?f?h?z?�? �?�?�?�?�?O
O,O RO@OvOdO�O�O�O�O �O�O�O__<_*_`_ N_�_r_�_�_�_�_����$SAF_DO_PULSڐ��o�84�a�PCANҚ��4�aF�"��"5�C��րր
@4a���ĵѵ�Xa�� ���o�o�o�o�o�o yo 2DVhc�o�r���rXaXad�x�q�q͑Tesy @�������y� �����_ �p.�T��.�k��}�����T D����ŏ׏����� 1�C�U�g�y����������ӟ�?�I��y���2�D�	���i�;׃oJ�i�p�l��
�t���Di��qhaJ�� � �g�i�ha`e Paӯ���	��-�?� Q�c�u���������Ͽ ����)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m���ߣߨ��+������� ��&�8�J�\��u ������������ �*�/�l�F�0)��� ����{����������� ����/ASe w������� +=Oas� ������// '/9/K/��o/�/�/�/ �/�/�/�/�/?|�5? G?Y?k?}?�?�?�?�?l0�����p��0%�0�0�0�d`q OO+O=OOO]GnO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o�o�g���d'���o ,>Pbt�� �������(��:�H�Q�~������q�w�M�	�12345678���h!B!S��e���pc  � ��$�6�H�Z�l� ~�������˟ݟ� ��%�7�I�[�m�� ������ǯح����� �1�C�U�g�y����� ����ӿ���	��گBH,�T�f�xϊ� �Ϯ������������,�>�P�b�t�߫;�j�ߪ߼������� ��(�:�L�^�p��`�������D��� ��� �2�D�V�h�z� ��������������
 ߯@Rdv�� �����* <N`r1��� ���//&/8/J/ \/n/�/�/�/�/�/� �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�?�OO&D߆AOSO`�/xO�O�O��CB��A��j   ���h2�b�} ��H
�G�  	ĩB29O _2_D_V_Rf\�ogL��1�@3 4 5 6f_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�oP�o�o�o�^P!r('r -?Qcu��� ������)�;�@M�_�q������A g@�h@Q�B<�� ���Q  ��ɋ㏖�ƂQQt�  �@����`��$SCR_GR�P 1"X��"al� � }��� �E�	 j��r���|�hA�������������䟬M���@�D�` D��@|]��'�ᛊ\�R-2000i�C/125L 5_67890PX�~PRC2L g����
V05.00 ������vS�H�B��r���a���a���S�������ǩ	��J�*�<�N�`�h���H�r���v��ѥh�D�y
��-�C3�����ݾ��B��r	��������XS�������¤@h��ፏh�  @��ȶD���?�XC2�r�_���%�ܟIϟ��;ϴEh�����B����B�  B�33BƘ��ŗ¨���A�@�����Ď�s@���� ?�����¾@
��ˎ�F@ F�`5�=�4�a� L߅�pߕ߻ߦ����� �����.��+�=�O�B�]��ߣ���� ��������!��E�0� i�T���{_���͟�������
����@+�&�,����R���h12#34f�x�F7O��A���������Y�$� �Q�� �'5JVh7  �����
/�"A�ECLVL ; !��Ѣ��"!L_DEFAU�LT*$}����uP>#HOT�STRJ-�"!MIPOWERF) ��EV%%WFDO�K& V%!"RVENT 11!1!w#� L!DUM�_EIP/�(�j�!AF_INExJ ?4!FT�/>>?b?!a�z?�;��Q?�?!RP?C_MAIN�?�8q��?�?�3VIS�?��9��?FO!TP&9@PU=O�)d5O�O�!
PMON_POROXY�O�&e�O��OYB�O�-f�O*_!�RDM_SRV�+_�)g_v_!RȊ�_�(he_�_!
��0M�O�,i�_o!?RLSYNw�*o�5g8�_Zo!R3OS�/�l�4Io�o�!
CE[@MTC�OM�o�&k�o�o!=	�bCONS�o�'�l�o>!�bWA'SRCE_�&m-�;!�bUSB��(ny�u?�9S�� #�H��l�3���W����'RVICE_K�L ?%�+ (�%SVCPRG1����2���3+�0��4S�X��5{����6�����7˟П򀃤��9� �_H���� p������E���� m��򁕟�򁽟8� ��`������5� ���^�ؿ��� �� ��(��֯P����x� �&����N����v� �������ƿ@�B� ���҂�ُ뀋��� ���������@�+� d�O�������� �����*��<�`�K� ��o����������� ��&J5nY� }������ 4XjU�y� �����/0//�T/Ɗ_DEV ~�*�MC:_/~q!GRP 2�%�� �bx 	_� 
 ,� 1@UK� p� � � U	� � \$�"��" =�$�!�  �$�%\#�#���!�!1P�!�!\+�#J� �$1577#\$�!Y99?  &8-5;C7
8]9�?�#�!%=�?��3�5�!1EO  Q � sa�1�!�%I�!�$+?0w� �� �!�+� 2>OGt� ]�� &� "� *� D�(�$�A�F!eI�5
A9� �$�9AO�# �!�5�?+[15%5t_�#�(O?;�!1�!q_ ?;	5=E�?C7�_"o1V�$s� �0�� �@�   %h-3�#D�q��H�8�?�#� A�D1mK?;Ua�8 =OkQ1�!�_S_1	O �oZA~ew�P�W���$�1�v4�o-��=�c�J� ��n��������ȏ� ���;�"�_�F�X���Z�}	�0X� ��D\!uu�  �� �Rd�a��C7�d�a1A � C7�a�!�o+��a�a�? W�}�����ʯ��� �@�$��H�/��u
T)�3�<�$Yk���U1��o��u�5�sG�5 ¯�.8%�?Ϙ!ə-5 ���W-ϗ�-9]����! տ_�A�>�9�b�I߆� ��߼ߣ�������� ��:�L�3�p�W��{� ����!��� ���$�� H�/�A�~�e������� �������� 2V =z���g�� �
�.@'dK �o�����/�/�</I)d �P�\6�� ����%�2!��A�� �}�M�9U��'l�I*g @x�A���3AiW�?�R�ZA��@�1���-������=u����=��%����o�-?,�@���8� @I	r?�3��@-vyI)%�PALLET_H�EIGHT_CH�EC�A? P��	�b%�����z������+�W�Bӝ�������V5�f!A�����o��A��v@� �@<��B���V=­|���� �.�7�Ң²����'V=�N�M>���9@0@��{�@�)RB�ZNV9%PL�ACE_4LEF�Tpb�? P���b%?;+��q��=@�+K;m�W~�F�V>U�n�V=�`�>��HFOB�C>�(��������CzV=B3+�A�������2S���*N�(�Ax������7?��q�@x;�?�߰��:�:R1�?�B,�P�&Wb%�R�����~�AJ� ������u��z�YV=@�w��&7�B,��V?�0����8@9�*N��W�������e:><-��_�e���Z�V=?����A?q���y��@/��@\4�?%��:�PICK_IN�COMING _�POIN�OW!(P�Ji6 ^B�s�B+=A��¾=\	A!�MB��>�������
Aߎ�#>�H@A��Aɗ�~>�
������>����?du´��B�7�5N^1��P?=b���h���%*��$�� ��v_�W�O�of$P���b%��b�������Eu�<d��,��B4ɴV=���;�� - �@�c5� �?�?�A����~>,��A
��<5�M��}iA����N^��@`a~���dpAK�����&p�м�p�?�;?�D�1�P�2f!:�m�u� ?�� ;������#|����>��{���:@��=;@�A��]zE�RN�(qAf,���vʷ�1j�ߜC"��N���/�`��B����>�-K����IA��zG�RIPPER_O�PEN ?ogPׯ��b ��"� ���f@H�=/�����ؽPl�>�����0A�&����ք�6�ߒ@ICmV=�4���������ƾ���w�$C#��N�����X%����?�o-?�?4�� �v|�Q?JACKPO�4叾�4P��66�#������E�������~fV>���d�7A��	 ?�4P?߿<BAt��~>��c��Q���\[W!¥
:B��8�>���^R��)�X��ښm@�'�B�<տ�;? D��)+663�~Bx���Bͼ��d�A���B��ɉV=>����J�AJ�*���P��+������RN��-�©�X��)ͱ °�/\B��>��Ԍ@p�b>��m�??a:,���iq��^�yg�-�7b%B*\A���s@oP�_��{AŁA���q�A�VAI�.A�%�A�ڼ@�G����bV>������@��>#��+��Q��B��ʦ>�G����K���f�r�g��&2���!��O�L��͔C��b%=?����t��>��}<���k�8�O<e��q�>p���G��A�Um�Oj{a�;@�S�XRO�E�A�������2P^"��V=�3`A+_�����@J��@�!�?������	FIND_TOTE OS,��T�;�<P�Z��b%��i�����@�S9�:�T�%�V������N��Q��vߋA��FA@5��@X4Pƾ����6��z�B�6��0������A�nq����0���>�?��.@��'��0�KB�T�f� ߜP�e<b%����m�l���\�ox:�W~��?�A�G٦>����j�JAh�.��v�Jﾌ��ƾ��+�?K�l�C�7Z����������.V>e]d�A^�A�'E��" (@�2�A
�����(���e�Zu=�i��-��-e-�����=P����z�{���D��a��b��:A9@�#��n��+�L���]���ڍ���h +=*��B�jz@�1��V�����������:;���ks����W��ؔ����hP=���<|Bf2Ij��"���A�q{�A���۸IA2���^�B�v���>�?�_�;h���¶���Mh��Np��������_�@&?'���0��ϴO���Бv�b �f!���X�A�$���ɝ�ꒈ��>�R�N�����h{Bv?h�0�7?�����*N�;\� �rb�<W�G����c�WC��V>FC�A��������@��Կ ����򙛃\���5P����b%A�a���H���.�f>���-��%x����z�"r�@���CA�����h@��A����~>�y����@%�`�2�,������N�m��bp{�%1�A� @�"�A�L�ߚ��;_̕��4b%:���@B��?�ъ�@?k�; BQN���h����A����o0���'<�� ƾ$@��B������~:�Y|>�!q��@���A���O���%��6s�	�3�P���eb%<��_?����6��2�?��<�圿�;@���AE�N�?�?����F�s~>���&@�/��O�����¤��B[[A��`�]�@V����^e?�8��!d��NMAIN I�C�5��3P��jR��e��߿z=ࡑ�g���o����N�=ք����A��f?k�)B��@D�Ŋb�����B��� ~�������,BUK�E��,@>�7���P���@�$F������;~��D�*��Zu�������@S�@M����z���N�{j��m���%���]M^!���#0f.4�PA�q�?�����r���+A�j�T�{B�E���B�������@v�A`ha�?0~3ѱ+���\s?' ����@���n@6�F����@��!�n�!��ۀ	�����;�Alk'��<�M��1�|A���������v����A�J��A�� ���4�B��B�Q@��	oQB�z�^O�>]�BA��&�a��Am��{��!�=���Ad�h=�^���~��?*��A�
����@Qž���E޿��������>6��^�j;I��R���nC|�=Ş�����X�L�;��3�>#:L�V_p �fXRž�V]���>���I����������~���i/A�Z}�Q��.�@$Y��f.�@�Akl �����rL�B�@��s0A���V��??V�@�$�I�2_�D_*o�1u�֖����BI�NB��9?�l>�����Ҭ�j�=�!��AG����,B�����@k�C	���s����.�?���»z���`�j�A'A���f��?��<�����҄�PATH�� �O � P��2R�l�U�?�{����:�<�@v ��	��r�2i����@�����$l@:R��@.�1Z���M�@)���A���@:�£�S�B��O�x�q�@Q���ֿ���ņ�R2s/�DÅ�/ �խ?���P��Bf �~�A������4��A�B?�>�W�r�����Aݖe@6Β��X����������]�u{��-_����C���j�(�>$����=�s=����z<�n0A����������Aa���)Pz>�)G����ĻY�3�>�5^;+N�rΎ`�����A��A>[p����p���������ܼ>�Aì�U����c}�^O����	�@�UU>�Z�m�#�@�fk�o����O�4�P��RŻS�rX ?u4�f¿DB�<0[=����T���&A�����@;�3�?7?��H�s��h���~ˡ��K@�^�r�����̌Z@�@?�������
��H�ֲ)��%���*�%?\�1�;п��Ž����r�*�����5A�`/?{��a@g%2:?����9�����~�V2��BBU�uj����������@V3h�y�݊�oT K ��r�]��F�G����J@�O�? (������?Wo�Z�	�����z�[ ����A��������b����Ĉ�dֿ)���iy�BV�{���%��)�BR3�BU����)`A*w!ҿpK��0�^%МD���E��j�A� �>|,����i���&���������'>�o"�S @1�ߝ?�rS���!��*�6��cD��X����BY�	Z�DK���_�"B����%�AO�d��A�ϸϝ�4��t���]������A��=������¥��)�zN������畱��A.�c?��:�^�*V�������ɾ����B��������f��ڞ���+����@?$	A�=Y�m|�/��(P���u�@Գ�3�9���� <J������b���7�~�c ���6A��>^�9�?ٿ�L@i�,f.��9��.�^���������±_��B|���P��A���:nA��j7�@�&p�?�l��G�$P���ݚF��/���ٻ?,X�������1�O?���JZ�<��3���������lk�����O�8B�����y@EV|���¥����^����k�B�NB"�.B+�~B���
� /.����5��� ������"�[7>8���is����b>���,:�30��c�xAd��?k�f.w�Aݟ�n�_��p��S�@�������G�B�l��A�>����@��zߌ��� �. ��5���������S��<�z��L��r�����B"����&v�Q,�^ґA+a�@�`�z� ⶏ�waw|���� ���^-����B�ܿ�.�t��=?%���
GRIPP�����P�
|��u;�f@(���>���s�	?h��;k$��^�����?�$AL�'���0�WSQ���yږb�WA5mߎ�~�&ʡ�ҿq��+UR~ΐ�d�n��~?������+{���[����/ �P��/�5>�4p�����BS@�?���V��?"��Z�Ì������v��A�z!A����@�m1V�z�+��� <�[����g������e9>@�����3�A�����4L��N��/���r*rDk�k=P���5��@`��`B��?�0�3{����6~?`AA�e?֑�A�NA�_��@S�XV�~p���a����|������F��`�+Z��|���� �B��������mv�Yy�F?X?=O|1�:�vaq@*l��;sx;���B	�>�E��Z�����h��A�2?R�Z忳P>w�����+�=�S��="¦���������J��C�c��������$'_f���V� `�TOP:`�/���"�I�u=����?���dS:�:T@'��=��D�ڞ	������A��?!����IӿH�boV΢$�@>�����8�a�ǤBL(<~��ę1�����/8��yL�D/���/�_S��Q����a<dc��E`�Aȣ<����[�w����^<��>@���@
���>��Af�@Sp6}��4��%?�����ɾu&|��NC"s�~���W���_�²C.t?�9��>���sJACK�PO�d�_�b%P���&��5yB�tEA𐽆�qA��3A���mv���J���A�6Z��1��_t��)�/.Z�v]���� �g���?��­>�C������A$�+&������\��
!'����Yr*	MID_POINT Pp�|:O�rP������w�O���`����A�;R*���A������<"�A����@b�:��ґ��3��tB7q�J�3@�V�)�"�
��o��A`a~�0�����$����H���_c��P��ö֫'��A]E�8������gA]�O�B,c�v�(��ukA�oq�?C`���^���Vξ����'�h7�Q������'�^�����@�-
��H���V��2*��j��_��W�P��VE��a���<�!?�9�yz��󲽧�C�Z��p� A��[Ӿ(��@��p@��r_����*��je��T��BL�=Fڞ�ꭿ����O�l>���J0�?��pr/�+�o��KVE���z�?��R߾tQ�;O�?R?!@���Z������8�A��h�?k�)��]M���p_B6)�A�уq���@��Jq�_�����ӻ޺�@��>?~�������A�Q������#���2=��I�u?���:�mW~�V�׼���q~������6@tT��-#�AD�v?�����۔�@������������@�C*|w~�^�8���B��A5d��?��@q�>���.���6��!�t�|�.?��[������߳��>����?}A����A��V@��^ٞN$��BV�פ��"Ж���M� �v��m	�v8GB��dA�'?�f������������VE?���?��ATx�<�A��b+h�?at�>5 ��-$A� l�������@�v /B�&��BI���v���-��!��"^%%A�x@0�0U�J�+@Z4^���᰺�V߁�,P��H�U�N�@���j�7����AcA=���q^@)����KjA�<�?��\	?���%:��4!���)�p�����qd�P�j`~�^?�%%���@�א?��PT2����x!�o�kS�/�9�P�#�]���9T�?^J���E��ś;�hx~>�K_����Z�����@����U�U��	�����v���Z,���>A��U�L���c���d�xB�������%B ��A^��CL�AMP_CLOS�E G �Q,���P�$�'	���()^?1YO���Ƣ�������>��b��d�7�;3�@�kq@�>o"���>����J��R�O���V�\C�����}�#��B����/��B"�@�������Z���P��A�*V7bA!�7���=h
�A=�������2��B�#$Z=/`�<�_������.����(7>�2���r�����L����A&����i	�������R;��\��;P��B�VE�@k�AO��@��)�>t$ @�@��ª�E:�2�>p�N�A�ec?����KA���>�������U�$.�	�r_���+B�s�vQ_�+@�Q����N�A��*HB
�Yz�$�}H�D��F�:����@@�������������\=��Sm���@? ���@A�0��O�ja���=�@��s��gQ�fC��>�`��~��B��Bf��~�KA��b�Xtȣ��K"V@�b����@�����[�c�@A�_e<����������A�0�������dy��`�>ꎽ=p��$o��>�>�4o��n�����O�>�{�A��AJ\!������!��3��\����	Ot�Ɵ�k��	��?�)�����Y?�H��X4P��%��A�7��@/�ߠ�Z�J���B�U�1������[Z��hBN��vN��/�G��?��k�]@�*@���@F��;����?�2�P��e�VE�1W���c�����y���:��HC?�RW5�J� B����pA����ܟ�?3J����C!���1����¾��{¤�O���O5A9�}�@�c��`�(нSv@>-����K�KHOM�E �?�OuP�i���be���#�T?*J=���:�R�`���J�b�,p�����A��<���?�0�7����� ��b����EZ����B�w��@���@75�����3A2�N@�.]Bl��?���_�j�r�j%=�p��A�����y�;
s	@�i�=Y�5B}����� �B���+�{�����/b�*�k���7�>3M$�q.���M����&A9D��������uX�?�%���f����סy�s}��������@��1��5�����t�
G���������6%�A��ؠA�A���j��������i�?�)���gK����`̮>�{B���8B�� ����M��%_��6�H�I ��P�x��f�p2���0�@ө)��G^��{w�i	�"�Q����V��:R��A�^��v��A��B��3��#*Y���?'� ����#��{����7�B�����TA�I����&8|DYt��F�J�@����@!>��<�?��HB��a�B�o���+�Aۀ	@A�Z}�J$l������ ������61?���T�5�C�����)b�@��S��&_'������&pA�+�Y�O �� @�J��c����?V�=v@p�<����k�1� �BY���v@.��@������ۦ@�!������z�MyB:,��@).���!Í��>����sB���A��;��kA�#./��ş�ı��"�̖�A��ۛ�*�����=A��&>��)�{��N
��B8. ?���N���?*Һ���� �D��e�4�xܛ������+f�PA����G߾@�~Ɓ�+��c
��N���5�P���ſK����9����p��߿p{ߜ=�v���,�^��A�-�@VrS>(���v���6�B�I�2��@���i�C�l��f����G������ڿ�V���. @��>#�8m� �P���A��Am��V��A� ���A�n�����@�=���������xA?(�@�:�@r��A��xy�����m�(������K�B��gh�^>�yK���?�P�����?�1���2�
~Z�TH�E�_CHECK|o��P��z���>6��AZ��?���!����>�?�b�����NϲA�G�?��X��&����"��v3���p�o�Kq@7~����h2]>����A�v��P��V����"���'��~_�<i���P�����F��A���?AI�����@�AzB�<��f������5A�ݞ?�����
��@��1�wʒ����?䞰��=��·�Q�����^>�~�>��s�F:�?�=����'f�������?�� P�����F�%�A��PAGʽ���g@흅B��Kf�����d�A��@�9����%����YN�!�B���aY��qǽ���±W`B�Ȁ^>�@p��b�8 >y����)��*�ck��	MID_�POI����h���P��)>5<��t����A���(��V��C�	����1����*��A��=��@�픊�R����+�*W(���6�1��[����-Ү�����^R��A���@)��@N1}�A.M�V������P�"�>5B����A���A(��}<J��A��z��$��n���J�*A�O��@��0&����.BsƁ��
]�?ݑa<��[·q!���b�ZN�v>����wɡ��O��#@����n�������Qe3���19��m�?e[J�������@m��=1��o�����[�A�I�@���qߍ���_R��>�2��NK�IS�ܾ�We��f��iQjj2<���@�ˡ���g��7�@V3�h@��JOG�Gja��<Qe:�~����?h���?v��E���>K/u<�c���.[�I��[�1A����3���P�&�R�����=���3����'�©x���R@ZN�Ԍ@��q��k������@$'f@���JR_SET�UPPROGRAYM��$�Nk~�;ň�� ��>\�: ��?�t��N^>0��c�9A�����Cz@�6Z�@�̿�&H�@���G������`���(��-��?�4����c�?���0�J0���ϱ����/�N��&&� �з=��b:"��Ӻ��(��-#��c0��A}���U��U@��S@���>�&E@�������+�����(��	��W�?�l����X?��d�n9,�ȥ��/��/�?�"�~�a����a�Q��-n�=���:+�D/=��`qx�A�Ň5�������D@E�uB?�E�@������9���=��(�;����B`@yT�Z�J@7xw?�?,4���E�?�9SG 3"�N�~���]@�s6�A D*��������Y�"�D�N�WSQ���5A�`@�p@��@��&�(��%�g���������u�"�&���:A��><�b?��&��j86�n0�fO�?]_�Qf	�6
��dc�T��6?D��#�,'�X����,�N���8������8XOA#����b>���!+������1r>@ş��U����-��z�2ө��B�o�� ��B�_@7]C/LAMP� ��3f�Qf�FJ��������[���< �+����Ү����YNA��V!�@��{@6Β�z�U�)�h[�������R�£�%���u��ޢL_��ɼ���^k<@����� ���y��(�,oHf�[�~u���l��ǟ�=��Ү������rA���?��T@"��?�2���^X�����J�>@����U�6���G^�>�,@A�(�u�^�����(����8_J[<� |Qg���$�A����A8l����؎A^�AD�L������M{A���=������r���J�ξl5|���\?�$B���^¶i�9��N��OA�+������?�.t�@`5Ͼ���Pv���>ϯ�!�p�
��
�m��>N���=ט <-��=�i=���h0�����A���?�Z�}�]zE�c��tl�ӆ�?��ѽuA��¶��:����>OA���~��@}�d=��>x�/����}�����Z���Va@��˧BX6���� �����&�yξ�
����?�<B��+0A�p�?��)&�3O��9��}����`��>¤�#���rN��=�h��pA.�@�1���:��:h�u�o�T�  %�p����jF����.�AsT�<O����W�3�N{�
�o��f��Af���A�A��@AZ}�4�(��6�p�[���g1���Z����^���E�����`�0U�#�����(�6^?� TES�P�g��ZŽQJ���dHG@0��:�W~�bP��Ϳ5�@u5�����A\�G��!��@�f��@p���,4��6P��ee��g�K�~�����G����3L?'E��w�e�r:"��B,��D�K�e���Z�=%����J@� �;τ�8�y����,B���]MA�*�����@Iӊ�)���.?P��⎾�n�����^��p������s^�����x?����e�����XA)"��A�%=�M��<[�4��bM�
�v��Z�A�,:�����<A��µ��y�{�@0L��.ߘ¹��Q�9����?�v@�7��P����@d6ſ�]����+���������^H`�w�=�&��i!��@(��^!~}@���A�ि�Oja@� A��P�Pr����>+����^��´Z��1g�������W��+�@�����F/�����w��HOME ԁ�z�u����T������z�Ԍ�_>9lZ�����;Z�^�a���D5�A���H��7�Q@���^�/3���}��]��d��A¬�}������$c*���&��-s�@N��q��;��%�V� !e_CH��qK���������*���+��=�J��~�������^[�	��E�5A�5����ݰ@����@��x�^�������������¨�+���7
��D'��/ �J\!@R����z<�����b�ER_OP�END�V�$�A��4;�����,�=XS��?�s�Q1��^G��@��A�L���h�@�y@��j�b8/����^��옾��\;¦������
��-$����e�i��@7;_̊2s�
� q�X�=���6}�A��iAKs����A-�>����F.�P����zA���@��+��C��@����B4����#g�;׾�r²Ǜ����
�i@�A#��g���H���7�@�+��sB������ϵ�Y:����@?�zA��7=������?���
����L�ڻ+A���b���@�߈�M�e
�C+��&�2���m� ��M��³�/��m.��I|@�J�3�Y�?�� v;�?����HT�  #P��j�ž�I@��� �E����V��Bb�>�!��
�����B�,�'@S��[��^�.��.�/�.ھi��L�<�����_$PJ[��nY@�0��"���9*��MAI PLAS�TICi��  �P�8<�~A����b�<�_`A��m=�.��ޮ����`@BJ���$��ڼ�/�@�����;�&��C��>0R��x(����I���yK�A��7������S���4����
����INC�OM�br?GE;P��I���2�t�@���d��~V�@U�<����Op�$�FA����?��r/�>��vޮ�����ø��l^�>@���W^q���b
�����A���=aj��٠���(\�8V"O4G&a_�R5B`a�$SE�RV_\0L  �:uHP�Aa2TOU�TPUA@?V�B`@2TRV �2���q�  (�"si�p��pb � 3�q]2TSA�V&``ZLYTOP1�0 2~Y d� � �� p � �J`2C`e� s�B`Ƃ�P��B`>*J`B`�P�qJ`��2c�d�*` 
�Vohozo�o�o�o�o �o�o�o
.@R dv������ ���*�<�N�`�r� ��������̏ޏ�����UYP�_NSFZN�_CFG y&�KSTmQ�U8�GoRP 2�F�Q� ,B   A����QD;� B����  B4S�RB21�VHELL;�
��V�PĒP\Y����RSR�����F�1�j� U���y��������ӯ ���0��T�e��Q�\��  �:a%@e�����s�s��Q*`1����޽����	`�Pm����HK 1��(bÿ`� �^{ύ϶ϱ������� ����F�A�S�eߎ���ߛ߭ߩ�OMM ����߬�FTOV_ENB=T:a�U�;�OW_REG_�UI�ORIMIO/FWDL���ޅ�^P�WAIT�ɐZ�x�XP<��Tu�T�IM<�����V�A<P��P�_UNI�T����YLC5�T�RY<��U�PM�B_HDDN 2~[ (`��a� W� x��s����������������$8�O�N_ALIAS y?)&iS( he�Q Zl~���V� ���);M_ q������ //%/7/I/�m// �/�/N/�/�/�/�/? �/3?E?W?i?{?&?�? �?�?�?�?�?OO/O AOSO�?wO�O�O�OXO �O�O�O__�O=_O_ a_s_�_0_�_�_�_�_ �_�_o'o9oKo�_\o �o�o�o�obo�o�o�o #�oGYk}� :������� 1�C�U� �y������� ��l����	��-�؏ Q�c�u�����D���ϟ �󟞟�)�;�M�_� 
���������˯v�� ��%�7��[�m�� ����N�ǿٿ����� !�3�E�W�i�ύϟ� �����π�����/� A���e�w߉ߛ�F߬� ��������+�=�O� a�s��������� ����'�9�K���o� ������P��������� ��5GYk}���$SMON_D�EFPROG �&����� &*SY�STEM*���@+ �RECA�LL ?}�	 �( �}3xco�py fr:\*�.* virt:�\tmpback�=>10.$2�02.21:19680 2;M_o}4a/p8��� }8�s:orderf?il.dat����J/\/n/}/mdb:�'/43/�/ �/�/{�&�/I? [?m?�?#?��?�? �?�/�/�/EOWOiO |/�/)O�/�O�O�O�/ �?�?0?A_S_e_x?�? _�?�_�_�_�?O�O ,O=oOoaotO�O!o�O �o�o�o�O_�_(_�o K]�o�_%8� �� oo�o�oG�Y� k�~o��o4�ŏ׏� �o��2C�U�g�z �����ӟ��
� ��.�?�Q�c�v���#� ����ϯ�����*� ;�M�_�r������:��˿ݿp�xyzr�ate 124 �������D�V�h�{�|�#�8:172�@"�4��������� ��@�ϳ�D�V�h�{�!���69.254.1�4&�4:16120 %�7���������tpdisc 0 �ߠҢߴ�E�W�i�|��tpconn 0�� �2�������z�:����=�O�a�t�1�����6�������~�5�͡�����K]��6��& :��p���� ��I[m���6 �������4E/ W/i/|//��/�/ �/��0A?S?e? x�%?��?�?�?� /�/,/=OOOaOt/�/�O�/<O�O�O�L�$�SNPX_ASG 2���Q��  �B%��O6_  ?���FPARAM �UQ ��	$[P9T� �9X�T�PPO�FT_KB_CF�G  �#U�CO�PIN_SIM + [�R�_�_�ocPRVNOR�DY_DO  �U�U#bQSTP/_DSB�^�Rgo��KSR Y� � & PN�S0001 PR�OGXQEIGHT�_CHECK�Y�sd�STOP_ON�_ERR0o�B�aP_TN Up��A�bRIN�G_PRM�oBbV�CNT_GP 2� U�QPx 	��V�YePs|}ZPr���p��t��w�JV}D7pRP 1!^Y�Pvqa���� �0�W�T�f�x����� ����ҏ�����,� >�P�b�t��������� ������(�:�L� ^�p���������ʯܯ � ��$�6�H�o�l� ~�������ƿؿ��� �5�2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ��� ����������*�<� N�`�������� ������&�M�J�\� n��������������� "4FXj| ������� 0BTfx�� �����//,/ >/e/b/t/�/�/�/�/��rPRG_COU�NT�V�r�)ENB�%M3�T?_UPD 1"�kT  
�/|Bd? v?�?�?�?�?�?�?�? OOAO<ONO`O�O�O �O�O�O�O�O�O__ &_8_a_\_n_�_�_�_ �_�_�_�_�_o9o4o FoXo�o|o�o�o�o�o �o�o0YT fx������ ��1�,�>�P�y�t� ��������Ώ��	�� �(�Q�L�^�p����� �����ܟ� �)�$� 6�H�q�l�~��������Ưد�����,_I�NFO 1#R5�80Z�	 �1�u�`�����<3��������������པ��������뾻����@k�፥����� D��z�?��C2����ݗ澹��DB�&�8�� YS�DEBUG� S0��(�d;9c�SP_PwASS�%B?u˿LOG $O��\1  (���?��(�.�  ��71(�
MC:\�Ģ��)��_MPC��� ����.����UD1��25��SAV %��1�l��*�Q�SVb��TEM_TIME� 1&��]0 �0 ��'���� 4�*�4�F�c4�p���MEMBOK  R571�����7�I�Y�X|�80� @Y�&��@{���t�������
��@���)�;� M���f�x����������� �����
.@@Rdv��,e� ����(: L^p�����`�� //��SK����!"�R/d/v/j��80  x/��/�62&�$����/�)(���!O�*�C=APC?_65>c�gⰆ?�d?�?�?�?���?�,��O9OKO]OoO�O(�$ �O�O��O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_�_o#o/�T1SVGUNS�PD�� 'u���F`2MODE_LIM '��y�Bd�2O`oa(��AeA�SK_OPTIO�Nj��y��a_D�I��ENB  ���u��aBC2_GRP 2)5%u��ј��@C�"s:lBCCFG +�kb(��2*�Yz`w �������	�� -��Q�<�u�`�r��� ��Ϗ���ޏ��'� M�8�q�\��������� ݟ���ڜ	�۟<�N� ɟ+���o�����̯ڪ 5%��������>� ,�b�P���t������� �ο��(��L�:� \ς�pϦϔ��ϸ��� ���� ��H�.��\� nߌߞ߰�.������� 
���.�@�R� �v�d� ������������ �<�*�`�N���r��� ����������& 68J�n�Z߼ ����4"D jX������ ��//./0/B/x/ f/�/�/�/�/�/�/�/ ??>?,?b?P?�?t? �?�?�?�?�?O�O .OLO^OpO�?�O�O�O �O�O�O __�O6_$_ Z_H_~_l_�_�_�_�_ �_�_�_ ooDo2oTo zoho�o�o�o�o�o�o �o�o
@.dO| ����N��� *��N�`�r�@����� ����ޏ̏����8� &�\�J���n������� ڟȟ���"��F�4� V�X�j�����įzܯ ���0���T�B�d� ��x�����ҿ����� ��>�,�N�P�bϘ� �ϼϪ��������� :�(�^�L߂�pߦߔ� �߸��� ���$�گ<� N�l�~������� ����� �2� �V�D� z�h������������� ��
@.dRt ������� *`N�:� ����n//$/�J/8/n/X&� �$T�BCSG_GRP� 2,X%��  ��  
 ?�  �/�/�/�/�*�� ?">�?E?/?i?{=�"�#.~�,d���1�?�!	 HC� {6&ff�2� {5Ƽ1A��!�?�9D;)�{6��F|4FAB4�?�?HL@�YA�8$B�:O�MCj���PN333{5B�C�O�O�O`{9�O_�N|4>�G&�AB�_Z]@�8[6 �8�U�_^_p_�_�_�_��_o#o2kh�La	�V3.002b	�rc2l2c	�*n`fd�"}o<fG�_?�33� X�a�i �`�m�o  ��# _�o�e�!J2ʗ#/�-�o
xCFoG 1X%�!��!4z��"�b4�x����z a �����+�� O�:�s�^�p�����͏ ���܏� �%�K�6� o�Z���~�����۟Ɵ ؟���5� �Y�k�q� �v�����D�ͯ��ݯ ��'��K�6�o��� ����`�ɿ���ؿ�� #ό!x/H�T/X�Z�l� �ϐ��ϴ�������� �D�2�h�Vߌ�z߰� ��������
���.�� R�@�v�d������ �������0���P� r�`������������� ��&8��HJ\ ������� �4"DFX�| ������
/0/ /T/B/x/f/�/�/�/ �/�/�/�/??>?,? b?P?r?�?B��?�?�? ~?O�?OO(O^OLO �OpO�O�O�O�O�O _ �O$__4_Z_l_~_8_ �_�_�_�_�_�_�_ o o0o2oDozoho�o�o �o�o�o�o�o
@ .dR�v��� ����*�<��?T� f�$�"�����̏���� ޏ ���J�\�n�,� ~�����ȟ������ "�ܟF�4�j�X�z��� ��į���֯���� �0�f�T���x����� ҿ������,��P� >�t�bτφϘ���H� ����
ߴ�:�(�J�p� ^ߔ߂߸ߦ����� � ���6�$�Z�H�j�� ���n��������� 2� �V�D�f���z��� ����������
 R@vd���� ���<*` rߊ�"�X�� /�&//6/\/J/�/ �/�/b/t/�/�/�/�/ "?4?F?X??|?j?�? �?�?�?�?�?�?OO BO0OROxOfO�O�O�O �O�O�O�O�O_>_,_ b_P_�_t_�_�_�_�_ �_o~�.o@o�_o ^opo�o�o�o�o�o�o $6HlZ| ~������ � �D�2�h�V�x�z��� ���ԏ
���.�� >�d�R���v�����П �������*��N�<� r�`�����Ro��ү� ����8�&�H�J�\� ������ȿڿ쿪�����4�"�X�B�  ~��� �Ɩς���$TBJOP_�GRP 22J���  K?���	�µ�4����R� ��� �,^��� �� � s � ���� @~���	 ߐC� 2�Qp�D������N҇&ffV�K�W�i�<�9]2�?���?L�͊�BH � A�Hץ߰�Ds)���>��SF�!Y����g��� �ҏ��>���<��~��?333?fh�~�B�  B ��<=���D5mF���n�w�ы��Af�����C+�&�.���Cj�����߁�����;ć�B�S��Ⴔ����]���������<;��6����F��� j�|�N�O��"(����z�J6���>_���C4(��� }������ ��&@*\f �r�������'/����ưJ!N�	�V3.00��orc2l��*t ���}��/�' F��  F�  G�X G7� G�R� Gr0 G��� G�@ G��� G�\ G��� G�` G��� H
� H�d H" H�.� H;� H�H2 HUޝ"E��� E� �!F�@ F� Fj` �F�� F� ��"�!� G$� G� GVص#��� G�L G��� G�h G��� =u=K+,XZ5����r?�2���3?� � &����ESTP�AR v�����H�R�0ABLE 15�� �0�0D)D����|:�'��(�(�ǉ��'	��(
�(�(A����(�(�(�6RDI�?���FA��@��7OIO[OmH�DO�O��K�O_ _2_D^�2S�O�� �Joo)o;o Mo_oqo�o�o�o�o�o �o�o%7I[ ���P�_��C�}�_�_ �_�_gOyO�O�O�O�H��2�rNUM  VJ���"���� @�@�2_CFGG 6k��&�@���IMEBF_TT��1����0��VER��CAÆ��R 1=7K 8/��3 ��P�
 M��  ���*�*�)�;� M�_�q���������˟ ݟ���\�7�I��� m��������ǯٯ�>��  PDT�&�� � "[L�^� �{!�M!�����UK���ѿ�_DE��� ��OTF,�>� �$1Cd�v� �$�������s�����RI�D���_e�چ@���0MI_CH�AN�� � ��D_BGLVL�����1��ETHERA�D ?�5�����00��:e��4�:71:d0:6k6 ��7��68�{69��ROUT׀!iZ!<�Z��9~��SNMASK������255.F��2.`#���5������0OOLOFS�_DI Tռ�O�RQCTRL !8��PS�?8�T'�\� n��������������� ��"4FXj|��K�����2PE�)�TAI����PG�L_CONFIG� >k�{����/cell/$C�ID$/grp1��M_q��KS� �����//� >/P/b/t/�/�/'/�/ �/�/�/??�/�/L? ^?p?�?�?�?5?�?�? �? OO$O�?HOZOlO ~O�O�O1OCO�O�O�O_ _2_�~}�Oh_z_ �_�_�_�_0���_�]��Oo1oCoUogoyo �O�o�o�o�o�o�o�o -?Qcu� �������)� ;�M�_�q�������� ˏݏ�����7�I� [�m���� ���ǟٟ ������3�E�W�i� {�����.�ïկ��� ����A�S�e�w��� ��*���ѿ������+�&�User View ;�}}1234567890\�nπϒ���϶Ͼ�G�����B�2Oɻ� �2�D�V� h�z�����I�3��� �������"��C���4��|��������5�����5k�0�B�T�@f�x��������6� ����,>��_��7��������Q��8�L^�p����� �lCameraM�C//0/B/T/f/DRE��/�/ �.Z��/�/�/??(?�  ���x?�? �?�?�?�?y/�?OO e?>OPObOtO�O�O�����/O�O�O__ ,_>_�?b_t_�_�O�_ �_�_�_�_o�O�Gj� �_Poboto�o�o�oQ_ �o�o�o=o(:L ^po�GD;	�� �����o<�N�`� ���������̏ޏ� ���s�(�:�L�^�p� ��)�����ʟ�� � �$�6�H�G�	ߟ ������ʯܯ�� $�6���Z�l�~����� ��[��G:K� ��$� 6�H�Z��~ϐϢ�� ��������� �ǿٷ9��a�s߅ߗߩ߻� b��������9�K�]�o���"	�0 ���������(��� L�^�p��������� �����������G Yk}��H��� �41CUg �[;����� �/�1/C/U/�y/ �/�/�/�/�/z���K j/?1?C?U?g?y? / �?�?�??�?�?	OO -O?O�/�%3k�?�O�O �O�O�O�O�?	__-_ xOQ_c_u_�_�_�_RO �%�{B_�_	oo-o?o Qo�Ouo�o�o�_�o�o �o�o�_�%��o cu����do� ��P)�;�M�_�q�<��*}  .y�� ď֏�����0�B��T�f�x�   C���o�2oD����?�-B�  C3�*q���ɺ�����*q@+� BS���h�[*p?�łBl@֑v������z�ǟ Aǒ^|"�\��x6FBo� Ο\�������̯ޯ� ��&�8�J�\�n��� ������ȿڿ���� "�4�F�X�j�|ώϠ�`��������&� 
*p�(  覀( 	 ��0��T�B� x�fߜߊ߬߮����ߠ����>�,��� ��������� ������%�,sr�O� a�s������������ ��8�'9��]o ��������� F#5GYk}� �����// 1/C/U/�y/�/�/� �/�/�/�/	??b/?? Q?c?�/�?�?�?�?�? �?(?:?O)O;O�?_O qO�O�O�O�O O�O�O _HO%_7_I_[_m__ �O�_�_�__�_�_o !o3oEo�_�_{o�o�o �_�o�o�o�odo ASe�o���� ��*��+�rO� a�s���������ߏ ��J�'�9�K�]�o� ��ȏ����ɟ���� �#�5�G���k�}��� ֟��ůׯ����T�4�@ /�<�N�`��/�6����)f�rh:\tpgl�\robots\r2000ic���_125l.xml�Ŀֿ�����`0�B�T�f�r���r� �ϩϻ��������� '�9�K�]�t�nߓߥ� �����������#�5� G�Y�p�j������ ��������1�C�U� l�f������������� ��	-?Qh�b ������� );Md^�� �����//%/ 7/I/`Z//�/�/�/ �/�/�/�/?!?3?E?tW>y��� 6����<< �� ?�W;�?W?�?�?�? �?�?O�?0ONO4OFO hO�O|O�O�O�O�O_��O�O_J_X��$�TPGL_OUT?PUT Ab�b�� z0��x6FB�PZR�ş�B4  �Qb���ɺ����ZR�5/�B�  �1��^��_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o%�7Ewz0�OPcel�l/cont1/�grp1/dcs�/cpcz/z6�/f �eB��?� �,kB�PX���q ��g�B^����X�7��@^���� ?�QBО�X��u:^��p�XO�r�u$[mx1y�u��p�q߼ZOBX��$9A�r�u��֊s<����v2345678901f�x����� ����ȃ�sd�����&�8�J��s}M�u��� ������U�g���� )�;�M��[������� ��˯c�ٯ��%�7� I����������ǿ ٿq���!�3�E�W� �eύϟϱ�����m� ���/�A�S�e��� sߛ߭߿�����{��� �+�=�O�a����� ������������'� 9�K�]�o�׍}u1��@����������
@|?�.@�: ( 	 Cuc��� �����;) _M�q���� �/�%//I/7/Y/@[/m/�/�/�/Qv�x0 �6�/?=�/5?G?!? k?}?Kz�/�?�?Z?�? �?�?�?,O>O�?BOtO O`O�O�O�O�O�OPO �O(_�O_^_p_J_�_ �__�_�_�_�_o$o �_0oZo�_�_�o�o<o �o�o�o�o ~oD V�oB�fx�� 2�
���@�R�,� v����p���Џj�� ����<���$�r��� ����������N�`� &�8�ҟD�n�H�Z��� �����쯆�د"�4� �X�j�ȯR���:��� ֿ�¿��|��T� f� ϊϜ�vϨ���0� B��ߴ�"�P�*�<� �ߘ��ϼ���hߺ�������:�L��")WGL1.XML
����$TPOFF_LIM � ��!����N_�SV��  ���P_MON MB�%�����2��STRTCHOK C�%�������VTCOMPA�T��H��VWVA/R D��k��� � �� �����_DEFP�ROG %��%  R_SETUP��RA�������_DISPLAY������INST_�MSK   ���INUSER�>���LCKGQUICKMENk���SCRE� ��%I�tpsc@��G� �	�� _�	�ST<���RACE_CFG E���k���	��
?��HNL 2F��� *r� ��^p �������ITEM 2GJ� �%$12345678901/C%  =<;/a/s/{#  !�/�+��E/�/��//�/S/? %?�/;?�/�/�?�/�? ?�?�?_?O?a?s?�? �?O�?gO�O�OO�O 'O9OKO�OoO_A_S_ �O__�O�O�O�_�_5_ �_ok_o�_�_jo�_ �o�_�o�oo�oCo�o yo9�oIo��o �	-�Q�#� 5��Y����e�}� �׏�M���q���L� ��g�ˏ�������%� 7� �[���+�Q�ן ǟٟ�����3�߯ ��{�;�����ï=� 篓���˿/�׿S�e� w���Iϭ�m��㿋� ����=���a�!�3� ��I߻�ߖ��ϱ�� ������]��ߓߥ� ���u������5� G�Y������O�a��� m����������C��y�+����xS�H}
�  �}
 "���
 ��+�
�UD1:\8����R_GRP �1I+� 	 @��� ������ $/�2*�8\/G/�/k%?�  �/�+�/�/�/ �/�/??%?'?9?o? ]?�?�?�?�?�?�?�?�O	K%O7O�S�CB 2J� �/�O�O�O�O�O�O��O__�UTOR?IAL K��^_�V_CONFIG L�z��_n\OUTP�UT M�	�P���_oo1oCo Uogoyo�o�o�o�o�o��o�Q�\Reg�ular Option�o0BT fx����������_�!�3�E�W� i�{�������ÏՏ� �d��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v������� ��п����*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x�����������������U� ���_9K]o�� ������� 5GYk}��� ����/1/C/ U/g/y/�/�/�/�/�/ �/�/	??,/??Q?c? u?�?�?�?�?�?�?�? OO(?;OMO_OqO�O �O�O�O�O�O�O__ $O7_I_[_m__�_�_ �_�_�_�_�_o!o2_ EoWoio{o�o�o�o�o �o�o�o.oAS ew������ ���*=�O�a�s� ��������͏ߏ�� �'�8�K�]�o����� ����ɟ۟����#��C�B�J�X��>�-��"\Re�gular Option����ί� ���(�:�L�^�p� ��5�������ѿ��� ��+�=�O�a�sυ� 6��ϻ��������� '�9�K�]�o߁ߒϥ� �����������#�5� G�Y�k�}��߳��� ��������1�C�U� g�y������������ ��	-?Qcu �������� );M_q�� �����//%/ 7/I/[/m//�/��/ �/�/�/�/?!?3?E? W?i?{?�?�/�?�?�? �?�?OO/OAOSOeO�wO�O�O�$TX_�SCREEN 1}NV�>��}��O�O�O__(_:_�O���Oz_�_ �_�_�_�_K_]_
oo .o@oRodo�_�o�_�o �o�o�o�o}o*�o N`r���1 ����&�8��\� ���������ȏڏQ� ��u�"�4�F�X�j�|� ����ğ֟���� ��0���T�f�x��������%�ү�$UAL�RM_MSG ?5�I��@ ʯ�: ��G�:�k�^����� �������ܿ� �1�~�SEV  ��c��ECFG� P�E�A � �5@�  A���   BȦ2Q��@�����l� �A �Qg����Gu4P���~���nP�3������ą�A�YxQ�e<'��TyQe��
��_Qf �$"��0QfL~��Y{Qf�:��X�Qf�!� ��NQf�o�GR�P 2Qy� 0�¦1	 2�����I_BBL_NO�TE Ry�T?��l�2�@�1����DEFP�RO�%� (�%CLEAR_�IO LOSE �CHECK T_ J�7:�l�W�%Ϝ�� ����������,�>��)�b���FKEYD?ATA 1S�I��Op �ǟ6�����������
��,(�=�4(POI�NT  ]EG � OON����tN?DIRECT���I�OICE`�TOUCHUP���� RE INF k�#`rY�}� ����/&//J/�1/n/�/����/�frh/gui/�whitehome.png�/�/�/��/�/?��&point�/<?N?`?r?�?6  �%look+2�3�?�?�?�? O��?�6indirec*?FOXOjO|O�O�>clos�$9O�O�O��O__0�&touchup6ON_`_�r_�_�_4�&arwrg5O�_�_�_o o�H5oGoYoko}o�o �o0o�o�o�o�o �oCUgy��, ����	��-�� Q�c�u�������:�Ϗ ����)���M�_� q����������%��� ��	��-�?�F�c�u� ��������L���� �)�;�ʯM�q����� ����˿Z����%� 7�I�ؿm�ϑϣϵ� ��V������!�3�E� W���{ߍߟ߱����� d�����/�A�S��� e���������r� ��+�=�O�a���� ����������n��� '9K]o����������+��� �4F�""�o��#,g/�_(O?INT  ]�� IRECT ��  ND�// CHOICE�|:/�UCHUPe/ f/�/�/�/�/�/�/? �/3??W?i?P?�?t?��?�?�?�?Ɲ&Ewh?itehom�D O�2ODOVOhOw�Fpoin�_�O�O�O�O�O��Oi/direc��O0_B_T_f_x__/in_�_�_�_�_�_<�_�AclosD�_�>oPoboto�o�Jtouchup�_�o�o��o�o�Narwrg�_@Rdv� �������*� <�N�`�r�����%��� ̏ޏ������8�J� \�n�����!���ȟڟ ����"���F�X�j� |�����/�į֯��� ���?��T�f�x��� ������ҿ����� ,ϻ�P�b�tφϘϪ� ��K�������(�:� ��^�p߂ߔߦ߸�G� ���� ��$�6�H��� l�~������U��� ��� �2�D���h�z� ����������c���
 .@R��v�� ���_�* <N`����� ��m//&/8/J/�\/3�j+�@ j/�/�/B�/�/�/ C�,�??�8OINT�  ]%?'? IR�ECT Q?R?  �NDf2}?? CH�OICE@?�?80UCHUP�?�?O%O OIO0OmOOfO�O�O �O�O�O�O�O!_3__�W_6��Uwhitehom&d�_�_�_�_x�_��fpoin/�o-o?oQoco�_i/direc
o�o�op�o�o�owo/in�o�!3EWi�oachoic�_������/touchup�.�@�R�d�|v��^arwrg ��ԏ�����.� @�R�d�v�������� П������*�<�N� `�r��������̯ޯ ����&�8�J�\�n� ����!���ȿڿ��� ϟ�4�F�X�j�|ώ� e_+����������� %�B�T�f�xߊߜ�+� ����������,�� P�b�t����9��� ������(���L�^� p���������G�����  $6��Zl~ ���C���  2D�hz�� ��Q��
//./ @/�d/v/�/�/�/�/ �/_/�/??*?<?N? �/r?�?�?�?�?�?����;�sP���OO'M�?IO[O5F,G_�O?_�O�O�O �O�O
_�O._@_'_d_ K_�_�_�_�_�_�_�_ �_o�_<o#o`oroYo �o}o�o�o���o &8JY?n��� ���i��"�4� F�X��|�������ď ֏e�����0�B�T� f�����������ҟ� s���,�>�P�b�� ��������ί�򯁯 �(�:�L�^�p����� ����ʿܿ�}��$� 6�H�Z�l�~�Ϣϴ� �������ϋ� �2�D� V�h�z�	ߞ߰����� ����
��o.�@�R�d� v��߬�������� ����<�N�`�r��� ��%��������� ��8J\n��� 3����"� FXj|��/� ���//0/�T/ f/x/�/�/�/=/�/�/ �/??,?�/P?b?t? �?�?�?�?K?�?�?O O(O:O�?^OpO�O�O �O�OGO�O�O __$_h6_H_�J[�����s_�_�]o_�_�_�V,�o�_�o  ooDoVo=ozoao�o �o�o�o�o�o
�o. RdK�o�� �����*�<�� `�r����������Oޏ ����&�8�J�ُn� ��������ȟW���� �"�4�F�՟j�|��� ����į֯e����� 0�B�T��x������� ��ҿa�����,�>� P�b��ϘϪϼ��� ��o���(�:�L�^� �ςߔߦ߸������� }��$�6�H�Z�l��� ����������y��  �2�D�V�h�z�Q��� ������������. @Rdv��� ����*<N `r����� �//�8/J/\/n/ �/�/!/�/�/�/�/�/ ?�/4?F?X?j?|?�? �?/?�?�?�?�?OO �?BOTOfOxO�O�O+O �O�O�O�O__,_�O P_b_t_�_�_�_9_�_ �_�_oo(o�_Lo^o@po�o�o�o�o���k���������o�o}�o);v, '�l��w��� ��� ��D�+�h� z�a�����ԏ���� ߏ��@�R�9�v�]� ������П����� *�9oN�`�r������� ��I�ޯ���&�8� ǯ\�n���������E� ڿ����"�4�F�տ j�|ώϠϲ���S��� ����0�B���f�x� �ߜ߮�����a���� �,�>�P���t��� �����]�����(� :�L�^���������� ����k� $6H Z��~����� ��� 2DVh o������� �/./@/R/d/v// �/�/�/�/�/�/�/? *?<?N?`?r?�??�? �?�?�?�?O�?&O8O JO\OnO�OO�O�O�O �O�O�O_�O4_F_X_ j_|_�__�_�_�_�_ �_o�_0oBoTofoxo �o�o+o�o�o�o�o �o>Pbt�� '������(��� *��� ���S�e�w�O�������,��܏�� �� $�6��Z�A�~���w� ����؟�џ���2� D�+�h�O���s���¯ ���ͯ
���@�R� d�v��������п� ����*Ϲ�N�`�r� �ϖϨ�7�������� �&ߵ�J�\�n߀ߒ� �߶�E��������"� 4���X�j�|���� A���������0�B� ��f�x���������O� ����,>��b t�����]� (:L�p� ����Y� // $/6/H/Z/1�~/�/�/ �/�/�/��/? ?2? D?V?h?�/�?�?�?�? �?�?u?
OO.O@ORO dO�?�O�O�O�O�O�O �O�O_*_<_N_`_r_ _�_�_�_�_�_�__ o&o8oJo\ono�oo �o�o�o�o�o�o�o" 4FXj|�� ������0�B� T�f�x��������ҏ ������,�>�P�b��t�����o ���>o ���ß՟ 睿�	����,�L� ��p�W�������ʯ�� � ��$��H�Z�A� ~�e�������ؿ���� � �2��V�=�zό� k/����������
�� .�@�R�d�v߈ߚ�)� �����������<� N�`�r���%���� ������&���J�\� n�������3������� ��"��FXj| ���A��� 0�Tfx�� �=���//,/ >/�b/t/�/�/�/�/ K/�/�/??(?:?�/ ^?p?�?�?�?�?�?�� �? OO$O6OHOO?lO ~O�O�O�O�O�OgO�O _ _2_D_V_�Oz_�_ �_�_�_�_c_�_
oo .o@oRodo�_�o�o�o �o�o�oqo*< N`�o����� ���&�8�J�\� n��������ȏڏ� {��"�4�F�X�j�|� �����ğ֟����� �0�B�T�f�x���������ү�����0�
���0���3�E�W�/�y���e�,wϼ�o��ǿ�� ��:�!�^�p�Wϔ�{� ���ϱ������$�� H�/�l�Sߐߢ߉��� �������? �2�D�V� h�z��������� ��
���.�@�R�d�v� ������������� ��*<N`r�� %����� 8J\n��!� ����/"/�F/ X/j/|/�/�///�/�/ �/�/??�/B?T?f? x?�?�?�?=?�?�?�? OO,O�?PObOtO�O �O�O9O�O�O�O__ (_:_�^_p_�_�_�_ �_�O�_�_ oo$o6o Ho�_lo~o�o�o�o�o Uo�o�o 2D�o hz�����c �
��.�@�R��v� ��������Џ_��� �*�<�N�`���� ����̟ޟm���&� 8�J�\�럀������� ȯگ�{��"�4�F� X�j���������Ŀֿ �w���0�B�T�f��x��$UI_IN�USER  ��������  y�}�_�MENHIST �1T�� � (��QP(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,181,1� �17 VERIFY�)�;�M�_���'���34,4� 1 ALIBR�ATION� EFT'�����d�v���7�TUPPRO�GRAM�ET,22 H��G�Y�������4��LAST�IC_PALLET_L��8���������Ϗ�148,2 � ��HEIGHT?_CHECK7�Q�0c�����53Э� 4���������)�����13��ACKPO��00 ��Ugy\|�,70FP��`��������� ��.@Rdv� ����� /�+/=/O/a/s/�/ /�/�/�/�/�/?? �/9?K?]?o?�?�?"? �?�?�?�?�?O�?5O GOYOkO}O�O�O0O�O �O�O�O__
C_U_ g_y_�_�_�_�O�_�_ �_	oo-o�_Qocouo �o�o�o:o�o�o�o );�o_q�� ��H����%� 7��[�m�������� ǏV�����!�3�E� 0_N�{�������ß՟ ؏����/�A�S�� w���������ѯ`�� ��+�=�O�a�𯅿 ������Ϳ߿n��� '�9�K�]��nϓϥ� ��������|��#�5� G�Y�k�V�ߡ߳��� ���������1�C�U� g�y���������� ��	���-�?�Q�c�u� ������������� ��);M_q�� $������7I[m�|���$UI_PANE�DATA 1V������  	�}c/�frh/cgtp�/flexdev�.stm?_wi�dth=0&_h�eight=10���ice=TP�&_lines=�15&_colu�mns=4�fo�nt=24&_p�age=whol�e��z�)prsimA/j/  }m/��/�/�/�/�/�/ ) �/?�/5??Y?k?R? �?v?�?�?�?�?�?O�OOCOz���� c@ �C�{$���2
%�3�@.1(%dou�b�@2MO+Hual��O
_qKitree �A_E_W_i_{_�O�_ �_�_�_�_�_o�_/o oSoeoLo�opo�o�ox�o�oVH � c@	 "��sO�O�OP3
&( �O�(%t#p3�o�khird��~/��� ��)��oM�4�q��� j�����ˏ��ݏ�� %��I�[�B���oq 	2W�.t ��ǟٟ����b�!� E��i�{�������ï *��ί����A�(� e�w�^�������ѿ�� ��ܿ�+��bB�� _�d�vψϚϬϾ�� ��U���*�<�N�`� �τߖ�}ߺߡ����� �����8��\�n�U� ��y����;�M���� "�4�F�X���|��Ϡ� ����������s�0 T;x�q�� ����,>% b�������� �E/(/��L/^/p/ �/�/�//�/�/�/ ? �/$??H?Z?A?~?e? �?�?�?�?�?�?o� ?/DOVOhOzO�O�O�? �O5/�O�O
__._@_ �Od_v_]_�_�_�_�_ �_�_�_o�_<oNo5o@roYo�o�oO-D��o@�o�o
.@)�o e�ET����� �R��3��,�i� P���t���Ï���Ώ����A��H+C%K��$UI_POST�YPE  +E�� 	 	�`�� �����Cs��QUICKMENw  �� �����_RESTOR�E 1W+E����*d�efault�K  INGLE板PRIM�m�omenupa�ge,1388,1,27N�������޼� m  d�290,1�����'��ʦB�T�f�x����� 4�����/��
�� .�@�R���vψϚϬ� ��a�������*�տ 7�I�[��ϖߨߺ��� �߁���&�8�J�\� �߀������s��� ����k�4�F�X�j�|� ������������� 0BT��	s� ������� >Pbt�)��������SCRE�?ǝuw1sc�u23$U33$43$53$63$�73$83!#TAT�~�� ֓+Ek�U�SER /,$ksT5#�$3�$4�$5�$�6�$7�$8�!s�N�DO_CFG iX����s�PDv!��)�No�ne��� _INF�O 1Y+EZ0Ԑ0%�u?�Hc?�? �?�?�?�?�?O�?4O OXOjOMO�O�O�O�O���G1OFFSET' \��^1�O� ��_'_9_K_x_o_ �_�_�_�__�_o�_ o>o5oGotoko}o�o �[ן�m�o�o
�o#��HUFRAM7��6D1RTOL_ABRTGB3_r�ENBhYxGRP� 1]�ӑCz  A��s�q1� �����(�:�[v���U�x1w{MSK'  �uZ1���[v�NDq%R9�%�AXIS_6_T���*�JR_EVN�gp��6�22^��K
 h1U�EVgp!td:�\event_u�ser\Џ+�C7�0� 0Fe�#�SP�)�.�spotw�eld`�!C6 ��f�x���d!�o?� ��2�ݗ���!��e� ��E�W�Я{������� ï<��`���S��� ��̿w�������8� ���n�ϒϤ�O�a���υ��ϩϻ� �WR�K 2_�)q8��b�t� Pߙ߫߆� ���߼�����;�M� (�q��^������ �����%� �6�[�m���$VARS_C�ONFI0`�K �FP��t�CCRG2c�J�O��ʙ�DA��BH�J�pC�J���*(?�: �$��M�R�r2i�K�l�0	q���@1�: SC130E�F2 *�� ����X��ș��50l1<A@C���' ����!NsIv��8�,0b�? B���� �Z�:/�;/&/ _/J/�/n/�/�//�/ �/�/�/%?�I?[?��TCC��j�z@�9h8���j ��GF���
�k�K �%�UF12 Aut�o �0 e se�t �R�� �h"u C
�1em�~�3456789012I�A� �0������H�������fX:���3��(.:$@8�@9� (?:�o=L�m ���y���%I��Ox��j����%�� �O��1��_%W[B -hOzO�O�O�_�O�H �_�__%_'_9_K_]_ o_�_no�_�_�o�_�_��oo#o5oGo~�1SOELEC넙���~�qVIA_WO:��l���p��,�		��`�o�G��P ǫp�iXqSI�ONTMOU� ���u��m�:���<t�1 �FR:\�s\D�ATA̟�0�� UD1:\ ��LOG�   �%��EX0�'� B@ ���s�D�iPend�ant 249 �.design.local;�[����= �� � n?6  �����p�ηt#`φ	  =������ 
 MC�vTRAINZ��2��dO�p����m��}��sOn�; ( 1[���
9������џ ���=�+�E�O�a��s�����z�ISSTAT o�9y� �=-2997.6�665: was� less th�an accep�table va�lue: -10�0.0)���$80_?SIDE_B4�g;_IS_GE�sp�;����
rpj ���\�HOMIN�pq/�E�����rq$q�aC$B�m\��JMPERR 2=r�;
  �o�� ���e���.�_�R�d� vψϚϬ�������ϰ�Dc�W�RE�ps\�|�LEXg�t����@1-eP�VMPHASE  ���j!r�OFFS_ET_ENB��u�OyP2�tu�F%��|���<cB�`A�1�`� ?s33���1cA��cEP��|��x��H��x��A���M�� �j ��5y���x<��t9�I�?��i� �����Ö0�������[�{3��1����E ��҅�&��Z��w ?�1����Ⱦ��{�1� ������!S���#�� ~������� + OAsh�� �����
/9 K]R/�'/�/�/ �/�/�]/�/5/*?<? k/]?�/i?�?�?�/�? �/�??OC?U?�?EO SOeO{O�?�O�?�?	O �O-O�O�O+_=_O_y_ �O	_{_�O�_�__	o s_o?o9o�_xo�_�o �_�o�_oKo�o�o�'5w[�TD_FI�LTE�yo� �f�t����o�� ������'�9� Ɓf�x����������ҏ����W�SHI�FTMENU 1-z�<�%�f� 1�D�j���z���ٟ�� �����W�.�@����d�v�ï��	L�IVE/SNAP���vsfliv܂�կ�b�IO�N ��U���menu����r���3��$���{b���MO���|n��zY�WA�ITDINEND�  ��Kᷲ�O9K����OUT�ูS,���TIML���W�G�y�Ϝ��+�|�J�|�i���REcLE������TM�������_ACT����u���_DAT�A }b�v�% � RIPPER_�OPEN���`�R�DIS1�-��$kXS��~b���p��J���Z�XVR���;�$ZAB�C_GRP 1�*���`,�h2���7ZIP���F�sc�o������z�MPC�F_G 1���� 0�o'���?�����`p�� �	�y�  <�T�  �=̫?���;�\ÿ���7�����غ������\���D��z�?��C2����5f��	����jv�
�e���&|��x�������������10������?��k^p|�f���b ����ݗ澹�D#B���
��o � �
 .X�����:.@5��ৰ�����_CYLINuDfq��� Јf ,(  */�.-�c/W/>/{/b- ��/�/�./�/g/ ???R?�/v?�?�? �/�?Y???�?�?O�?`m?NO`O�?�2���x� ���O�o���O�_\�O8_�g��RQA��SPHE_RE 2��̲? �_O�_�_�_�_0OC_ o0o�?To�_�_�oqo �o�oo�o�o=oOo, �oP7I��o��l�9�ZZ�� ǳ�