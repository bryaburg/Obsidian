��   �A��*SYST�EM*��V9.1�0170 9/�18/2019 A 	  ����HAPTIC�_T   8 �$ENABLE�  $BBLNOTEENB=�MAX_ALAR�MSLIO=  ݟ&ALM- � $ERRCsOD<' STY;� 1&IO- �X �
$IOT�YP<$IND�EX�TRG�R�SRV1�VAL�=�2�3=�H�PCFG- $� 6$DEB�UG=COMP_�SW=	 �$$�CLASS  O���C��f���f8VERSIO�N@  �Z��* / a�f��l�
ܒr_DF� 2�C�( �  � #j�5���C��D�2 ������/./ @/R/d/v/�/�/�/�/��/�/��F�   D`�<	"�9G��CG��;2
84`8@9x?�?�?��?�?�?�?�?�d 2?6�
 +O=OOOaO sO�O�O�O�O�O�O�O$_�+Uu >
	/K_]S�3U��_�_�_��_�%P_MOT_	C��R