��   �A��*SYST�EM*��V9.1�0170 9/�18/2019 A 	  ����HAPTIC�_T   8 �$ENABLE�  $BBLNOTEENB=�MAX_ALARMSLIO=��&�ALM-  �$ERRCOD�<' STY; 1�&IO- X ��
$IOTYP�<$INDEX��TRG�RSR;V1�VAL=��2�3=�HPC�FG- $ �6$DEBUG�=COMP_SW�=	 �$$CL�ASS  �S��C��f��f8VERSION@�  ��Z��* / a#f��l�
�r�_DF� 2C��(  � � #�5Z���C�D�q2 ������/./@/R/ d/v/�/�/�/�/�/�/4��F�   `�Q<	"�9G���CG��;284`8@9x?�?�?�?�? �?�?�?�d 2?6�
 +O=OOOaOsO�O �O�O�O�O�O�O_�+�Uu >
	/K_]S �3U��_�_�_�_�%?P_MOT_	C��R