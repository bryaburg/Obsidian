��   �A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����FSAC_L�ST_T   �8 $CLNT�_NAME �!$IP_ADD�RESSB $A�CCN _LVL  $APPP � X�$8 A~O  ���z�����o VER�SIONw�  �Z�$'DEF\ w { ��� ���ENOABLEw ������LIST 1� �  @�!�������
[.@�d� ����/�3// W/*/</�/`/�/�/�/ �/�/�/�/??S?&? 8?J?�?n?�?�?�?�? �?O�?�?OO"OsOFO �OjO|O�O�O�O�O_ �O�O6__\_B_�_f_ x_�_�_�_�W