��   ��A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_  �$$�CLASS  O�����D���DVERSIO�N  ��Z�8LOO�R G��DD<Z$?���q���M,  1 <DYX< [�����D'�i�����iO/a/s/�A/�/�/�/$ ��/�/�/	;�$MN�U>A>"�� � <i#E?  �ı� ę� Ę ��0=?O?�5��s0Ĝ� ė����4y?�?�5D�
�0�k0���x?�?`7߰� D��0�@ذ?�?<J��'��P�5,O>O�:D�1�Z@ �?/�O���O�O�O�G�:�P�ݺu����T:u��g%P�9���:�O=� Y&�%P�DɸdC�?���QS��P%Pj����;��J:����%Pr�{�껁��Q;|�%P �Ħ
��Ķ���ZUU�I/�_�U�A;/#Q�����\�;Go�;��g�?����,��D0<�-a?�D��{��������Q7NUM�  ���a�� UfC2TOO�L%?\ 
;8^����w�z�̉��h�^��<.�����*��Z����C���,�x�Dj>>�I�� �]�׮Q�a?� ���.3���4�;�/��XC���m�a�i4 :�f3	o9�iD �mO�_'U; �_�q����� 	���?�%�Gu�[��4dc[!j	��