��   ��A��*SYST�EM*��V9.1�0170 9/�18/2019 A 	  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41�� d =R��&J_�  4 $:(F3IDX���_ICI���MIX_BG-<y
_NAMc gMODc_USd~�IFY_TI�w ��MKR-�  $LI�Nc   "_SIZcg�� ��. X $USE_FLC 3!p�:&iF*SIMA�7#QC#QBn'SC�AN�AX�+IN��*I��_COUN�rRO( ��!_TMR_VA�g#h>�ia �'�` ����1�+W[AR�$�H�!��#N3CH�P�E�$O�!PR�'I�oq6�OoATH�- P $E�NABL+��0BT���$$C�LASS  �����1��5��5��0VERS��7�  �Z��6/ �55�������@MF!�0�1RE��%�1{O��wO�O����#EI2.K!�O_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_oo�O+ �W?H9@ ���\j�0lo~o�i�ܧ � 2.I  4%BG���o���aP�|H%�o�g_A�oA  ewV���� �����=��.�@�c$"+ �kdK@����RA��X�� �1@fNʏ܏� �� $�6�H�Z�l�~����� ��RF_A��_A֟��� ��0�B�T�f�x���@�������4JM4��c6C!2�l��� /�A�S�e�w������� ��ѿ������(�:� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~ߐߢߴ������� ����2�D�V�h�z� ������������
� �'�@�R�d�v����� ����������#� <N`r���� ���&1J \n������ ��/"/-?X/j/ |/�/�/�/�/�/�/�/ ??0?3h�4�0v�g? @