��   ��A��*SYST�EM*��V9.1�0170 9/�18/2019 A   ����DCSS_C�PC_T  �4 $COMM�ENT $�ENABLE � $MODJG�RP_NUMKL�\  $U�FRM\] _VT�X M �   �$Y�Z1K �$Z2�STOP�_TYPKDSB�IO�IDXKE�NBL_CALM�D�USE_PR�EDIC? �EL�AY_TIMJS�PEED_CTR�LKOVR_LI�M? p D� L�0��UTOOi��O^*+&S. � 8J\TC�u
!���p\� E&|Y0  � �CHG_SIZ�O$AP!�E�DIS�]$!�!C_+{#s%O#J�p 	]$Jd#� �&s"�"�{#�)�$�'�_SE�EXPAN#N��  ,$STAT�/ DFP_�BASE 5$0K$4!� .6�_V7>H73��&J>- � }�n\AXS\UP��LW�7������d4r � < w?�?�?��?�?��//	0&ELE}M/ T �&B.2NO�G]@%CN�HA�DF#� $DATA)a6e0 � PJ�@ �2 
&P5� �� 1U*n   _VSiSZbRj0RjR(�VyT(�R%S�{TROBOT�X�SARo�U�V$C�UR_��R DSE�TU4"	 �bAI�SP_MGN�I?NP_ASSe#� PB!� `CiH�77`e��.fXc1�CONFIG_CHK`E�_PO* }dSHR�ST�gM^#/eOT�HERRBT�j_G]�R�dTv �ku,�chT1r
0R HpLH�d� 0  lt<xNe'AVRFYhH�^t�5�1� ��W��_A$R�4S;PH/ (G%�Q�Q�Q3wB;OX/ 8�@F!��F!�G �r{�zT�UIRi@  �,�F�pER%@2� $�p -L�_SF��D(��ZN/ 0 �IF(@�p��Z_��0�_�0wu0 � @�Q7yv	
�� _�$$CL` �2�����Q��Q��V�ERSION���  �Z��$' 2 �Q�  C�ell Box �In��*�h� ���m�����E�"� œ�����E� ŷ�����?Ĩ� D�ğ�����  d����Cz  ����:����JackpotT�Out_�q�w�,�����c��@���?�^� DH��Κ�@ȯ+���9�'��I�Incomi�ng[�n�����a � E	����D\ G �ȩ���ޡ�ÿ -���;�)�G�H�l� {���oϬ�������h����%�7�I�MiddleT�h�~���?9  �8`L߫�?C�&få��Οl�
��`15���C��1�G�Left Side�`�u��ߐ�O;� E�߭�CԐ�����Д�  D���������D�B�>D�Righg�z� �������ྱ���� ��Q��%�K�9O��ICK SLOW�DOW�z�߃�"ؐ�������ě����n�0BW�b�d�J2 SlowdowZ�������������[�C ې����1/E/_�h�z����D�����/ #/5/?I?Sπ?wω� ���?�?�?�??1? C?U?g?|O�O�?�?�O �?�O�O�OO-O?OQO�f_Y�pick d?cs tesb��)d����_��Ö@P�P�_`��ې�Qo_ ._@_R_TorO�o�O�O �O�o�o�o	o*o<o No`oro���o�o� �o���&8J\ ������p��̏ ��"�4�F�l�j�|� �����ďٟ���� �0�B�T�f�{����� ����������,� >�P�v�d��������� ί����(�:�L� ^�p��ϔ��ϸ�ʿ�� ���'�6�H�Z� � nߐϥߴ��������� �#�2�D�V�h�zߏ� �߳����������� 1�@�R�d�v�x���� ���������-<� N�`�r��������� ���)�J\ n�;����� ��%/7/FXj� ���/@/���// !?3?B/T/f/x/�/�? �/�?�/�/�??	O/O AOP?b?t?�?�O�?�O �?�?�?_O+_=_LO ^OpO�O�O�_�O�_�O �Oo_'o9oKoZ_l_ ~_$o�o�_�o�_�_�_  o5GVohozo�o �o��o��o�o� 1�C�U�dv���� �ӏ��*��
�?��Q�`�r�����������$DCSS_CS�C 2��ۑ�Q  P�100% S�afe Spee�}�b�l�F@
�,�ł�j�di1��j�C���'�,�
����i�����d�����ԯ 5���Y��i���R��� v�׿��������1� U��y�<ϝ�`��τ� ���Ϻ����?��c� &߇�J�\߽߀��ߤ� ���)���9�_�"���F��j����ΔGR�P 2ۛ ��ÄC��\En�њC  E5�� 	��5�ǀ#� \�G���k��������� ������F1j U�y����� �0T?xc ������/� />/)/b/M/�/�/�/ u/�/�/�/�/?(?? L?7?p?�?�?_?�?�? �?�? O�?�?6O!OZO lO~OIO�O�O�O�O�O �O_ __D_V_h_3_ �_w_�_�_�_�_�_�_��_.oŝGSTAT� 2ۙ-��<� ��?]����� 9�EL������]�����2F;���;˛f��2�D�J�O��ODIۑ`<jf�;����Ɓ�2%=g4�t�?�  �a��`4���ZC��@���Ɓۑje����S<��?t��M�tg�<￾�����i��Ʉ@>F �D��Yx�i>G[����0?}�}�<���a���Ϳ}��<����>W�A�,�]�9v�D�9�]{F�+�So?}�)BsÊJq�� ����.��ϳD�.��UzD~ܫ��i?���?�;~�=p�p�.;ϵ����?��˙?�b� no�o�o�gە�0�ە �\�n�H��������j �`iҏk�z���� 	�+�-�?�a���u��� ş����ߟះ�=�O� ��[���_�q���ͯÏ ���%��-��%�G� u�[�}��������ǿ ٿ��)�+�ѯkϝ�W���ϳύ�������?]��`�  �9��q�pq�]�������;�X7�;˒��p1�`��OγDI���o�3��"�b2%T��`�bS��`}3�d;�	+�o��<�#�`W��`�<�߸pN�f���t >F�@p~{J���u2p]<�"�N�>p6Bp�<����>[YA�6_��9��Vp_{�ټ+��np	����G�ѽ"��p&�ϧ��p��U&dD~�)��|�'C;}綬=�p&;���5��Vٻ��.�p1�(�
��.� �Ϻ������������ 8�J��2�t�Fό��� ������������( @^DVx�L�� ���0
Tf \�������� �/�/D/*/</^/ �/r/�/�/�/n?6 �/:?L?&?p?�?\?z� ��2�D�V�h�zߌߞ� ����������
��.� @�R��O�?�?�?d?V_ h_^?t_�_x_�_�_�_ ��/o�/(oFo,o>o `o�oto�o�o�o�o�o �o�oB�/r��_ p������_F ,�Z$�F�t�Z�|��� ������Ə؏��(�� 0�^�D�
������֟ �����_(_�? �?�?OO(O:OLO^O pO�O�O�O�O�O�O�O `�B�T�f� ����� �:��&�pς��j� ��~�����������*� �2�`�F�xߖ�|ߎ� ���߄�� �R��V� h�B���������� ��������F�,�N� |�b�t����������� ����<n�(r�^ �����Ŀj�|��� ����į֯����� 0�B�T�f�x����� ���/�/��/�/ �/�/??��H? `?~?d?v?�?�?�?�? �?�?O2OO*OLOzO  �O�O�/�O�O_�O (_:_0?~Od_�O\_~_ �_�_�_�_�_�_o�_ o2o`oFoho�o|oB_ �o
_�o �oDV 0N/`/*<N `r������ �//&/��z�� 8*�<�2H�r�L�^� ����T_�o䟶o���  ��4�b�H�j���~� ��ί��Ư���oF� X���D�����z�Ŀֿ ̟� �.����H�.� P�~�dφϴϚϬ��� �����2��޿tߦ� `ߪ߼ߖ�������� ���������  �2�D�V�h�z����� ��4��(�:����� ����������DV �>߀Rߘ��� ���4Lj Pb��X���& �*/<//`/r/h� �/��/�/�/�/�/?  ?"?P?6?H?j?�?~? �?�?�?z/OB/�?FO XO2O|O�OhO����>� P�b�t������� ������(�:�L�^� �_�O�O�OpObotojO �o�o�o�o�o�o�/�? �?4R8Jl� ��������  �N��?~����o|�Ə ؏�����R�8�f� 0�R���f��������� �ҟ��4��<�j� P����ޏ�����ί��*�8��$DCS�S_JPC 2�"�Q (� DRigh�t Side C�lear����C_9  @@��
#P}"QLefn��������Õ�����In j�����V��C*�� ����C򰮶����!��/"�`{�B�����At Pi�ck���A  ����$�
RH J?ackpot�����C!���L�߇��a�ݳkό�Sߡ������Home J1���˿ٙ���ff4���2���?�����������3������G��3_�G���4a����������5����¤  �ɤ����6������>���at� EOAT ch�g ���B�ffB�R�f��/�?@Fff@�����_�s��������������&` ?��vߨ�����b j���d��+�?�B� � B�bdsbl�� f����� �������2�������.�3J��
�'�{4���"Q�t����5 a�L�� �j��6��� B�>/�ߥ/�����F�2 limYiO�.�B�
�P����#��/�/?#P �/m?�/�?`?�?�?�? �?�?�?�?3OOAO&O {OJO�OnO�O�O�O�O _�O�OA__"_4_�_�X_�_|_�_�_�_J�S�S�W�L  a�fe Speed,�_»Bȉ�H񋤄1aG�2&`to�o7�A8��aaai��ro�o�_ �ofa�o�o?c *�N�r��� ���;�M��q�8� ��\�����ݏ���ȏ %��3��m�4�F�X� j�ǟ��럲��֟3� ��W��{�B���f�x� ���������A�� e�,���P���t�ѿ�� ߿�������s� :ϗ�^ϻς��Ϧ�� ��'���K��$�6ߓ� ��l��ߐ��ߴ���� 5���Y� �}�D��h� ����������C� 
�g�.���R���v��� ����������?Q u<�`���� �)�7q8 J\n����d�MODEL 2>kx^!���$<�c�X �B�fÈ  �A`  CHp �ǀ �o$F/X/�	zp xp$6  ë$�/�/j&�t(� �/�/@�&�!�%�#�9�! �hM7b?9?K?�?o?�? �?�?�?�?O�?�?LO�#O5OGO�WJ3 4�O=-=C\�(s ��s ��� �@CW �CbOtO�O\O__e_ <_N_�_r_�_�_�_�_ �_o�_oOo&o8oWo�\ono�o�o�o�o��L�o�o\�oE Wi{����� ����/�A���e� w�ď������я��� B��+�x�%S�e� ҟM���͟���P� '�9���]�o���ί�� ���ۯ�:��#�5� ��Y�k�������� ����ۿ�ÿ1�Cϐ� g�y��ϝϯ������� ��D��-�z�Q�c�u� �ߙ߫�������.�� �)�����#�Q�c�9� ��������<��%� 7�I�[�m��������� ��������!nE W�{��u���� ��F/|Se �������0/ //f/=/O/a/�/�/ �/�/�/�/?�/?? �t?=?O?�?�?�? �?�?�?�?�?O#OpO GOYO�O}O�O�O�O�O �O$_�O_Z_1_C_U_ g_y_�_a?�_�?�_�_ 2o	ooho?oQocouo �o�o�o�o�o�o );M�q�� �������_`� �_)�;������ޏ�� Ǐُ&����\�3�E� ��i�{���ڟ��ß� ���F��/�A���e� w�M�_�q�������� ��+�=�O���s��� ҿ����Ϳ߿��P� '�9φ�]�oρϓϥ� �������:�կ�� 'ߔ��}ߏߡ߳��� �����H��1�C�U� g�y����������� ��	��-�z�Q�c��� K�]ߋ���
���� R);�_q�� ����<% rI[m���� ��&/������/%/ �i/{/�/�/�/�/�/ �/�/??/?|?S?e? �?�?�?�?�?�?�?0O OOfO=OOOaO7/�O [/�O�OqO�O�O>__ '_t_K_]_o_�_�_�_ �_�_�_(o�_o#o5o GoYo�o}o�o�o�o�o �o�O6�O�o~U g������� 2�	��h�?�Q���u� ����揽�Ϗ����R�)�;�M�f��$D�CSS_PSTA�T ������Q   �t���ɐПԐ � Ν (�g  �x����͚��ԟ;�� W� t���k�損�����e�����¯p����鮦�SETUPw 	��B�x� k���4���U�D�y��h�����T1SC �2
�f�m�Cz�k�ݿ�ͺ�CP [RȼD�D. L�^� �ϔϦ�u��� ���Ͻ��$�6��Z� l�;�}ߢߴ߃����� ���� �2�D��h�z� ��[���������
� ��.�@�R�!�v����� i����������� <N`h�8ύ�& ����/� SewF���� ���/+/=//a/ s/�/T/�/�/�/�/�/ ?�/�/9?K??o?�? �?b?�?�?�?�?�?O #O�?GOYO(O}O�O�O p�O�O�OpO__1_  _U_g_y_H_�_�_~_ �_�_�_�_o-o?oo couo�oVo�o�o�o�o �o�o);Mq ��d����� ���I�[�*���� ��r�Ǐُ돺O�!� 3���W�i�{�J����� ��՟���ȟ�/�A� �e�w���X������� �����֯+�=�O�� s�����f���Ϳ߿�� ���9�K�]�,ρ� �ϥ�t������ϼ�� #�5��Y�k���Lߡ� �߂����������1� C��g�y��Z���� ������	���-�?�Q�  �u�����h������� ����;M_. ���v���� %�I[m<ߑ ��<����!/ 3/E//i/{/J/\/�/ �/�/�/�/?�//?A? S?"?w?�?�?j?�?�? �?�?OO�?=OOOaO 0O�O�O�OxO�O�O�O �O_'_�OK_]_o_>_ �_�_�_��_�_�_�_ #o5oGooko}oLo�o �o�o�o�o�o�o1 CU$y�Zl� ���	���?�Q� c�2�������z�Ϗ� ����)���M�_�q� @���������ݟ�� �_%�7����m��N� ����ǯ������ޯ 3�E�W�&�{���\��� ÿտ�������A� S�e�4ωϛ�j�|��� �ϲ���+���O�a� s�Bߗߩ߻ߊ���������'�9���$D�CSS_TCPM�AP  ����g�Q W@ ����w������	�
��������  �������R�����U����U �!�"�#�U$�%�&�'�U(�)�*�+�U,�-�.�/�U0�1�2�3�U4�5�6�7�U8�9�:�;�U<�=�>�?��@W�UIRO 2]g��x��� ������������  2DVhz����������� 3EWi{��� ����////A/ S/e/��/�/�/�/ �/�/??+?=?O?a? s?�?�?�?�?�?�?�? |/O�/9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_O�_�S�UIZN 2.g�	 �x�v��_ �_o��_4oFoXoo |o�o�ooo�o�o�o�o 0�oTfx; �������� �>�P��t������� m�Ώ������(�:� ��^�p���Q�����ʟ ��� ���6�H�Z� �/�����q�Ưد���_Z�UFRM R.f����8�@� R��v���c������� ���Ͽ�*��N�`� ;τϖ�qϺ��ϧ��� ��+�8�J���n߀� [ߤ߶ߑ�������� "���F�X�3�i��� {���������#�0� B���f�x�S������� ��������,P b=��s��� ��(:�^p K������� /$/�H/Z/5/~/�/ k/�/�/�/�/�/
? 2?D??h?z?U?�?�? �?�?�?�?
OO�?@O RO-OvO�OcO�O�O�O �O�O??*_<_�O`_ r_M_�_�_�_�_�_�_ oo�_8oJo%ono�o [o�o�o�o�o�o�o_ "4�oXjE�� {������� B�T�/�x���e����� ������,�ˏP� b�=�����s���Ο�� �����:�L�'�p� ��]�������ܯ�ȧ