��  	��A��*SYST�EM*��V9.1�0170 9/�18/2019 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP�fBI�IZ@� LRM_REC�O"  � AL]M�"ENB���&sON�!� MDG/� 0 $DEBUG1A�"d�$�3AO� ."��!_�IF� |� E/NABL@C#� �P dC#U5K�!M�A�B �"�
� O�G�f 0CURR�_D1P $Q3LIN�@S1I4$D���APPINFOE�Q/ �L A� ?1~5/ H� �79EQU�IP 2�0N�AM� ��2_O�VR�$VER�SI� ���~0C�OUPLE,  � $�!PPV1C'ES0�!H1�!"�PR0�2	 � �$SOFT�T�_IDBTOTA/L_EQ� Q1Q@�NOTBU SPI_OINDE]iEXBSCREEN_�4�BSIG�0�OKK@PK_FI�0	$THK�Y�GPANE\D �� DUMMY1�d�D�!�E4�A���ARG1R�
� � $TIT1d ��� +Td+TP� +TP+T5)V6)VU7)V8)V9)W0)W�2W�A+UFW
Q+UZW1
dW1nW1xW 4V�R~�!SBN_CF�![�0$!J� �; 
2�1_CMNT��$FLAGS�]�CHE"$Bb_OPT�2�� �ELLSETUP�  `�0HO��0 PRZ1%ocM�ACRO{bREP	R�hD0D+h@��bl{�eHM MN�yB
1�0UTOB �U�0 �9DEVIC(ST	I�0�� D@13�r�`BEdf"VAL�#ISP_UNI��p_DOv7=yFR_F�@K%D13�x/A�c�C_WA3t��awzOFF_�0N.�DEL�xLF0q8�A�q�b?q�pF�C?�`�A�E�C#��s�ATB�t�1�MyO� �sE � �[M�s��&�RE�V�BIL:�!X�I� �R  �� ODq`^��$NO`M�!QV�l�/�"i��� w����!X�@D�d p E R�D_EV��$F�SSB�&K`KBD�_SE&uAG� G
�2 "_��B�� V�t:5`ˁECY`�a�_EDu � �S C2�}`S�p��4%$l �t$O�P�@EB�qm�_O�KԂUS�1P_C�� m��d\�U �`LACI�!�a����� �:qCOMM� �0$D��Ñt@�pL��O��B BIGALL;OW� (KD2:�2�@VAR)�d!|AB �`BLO@S �� ,K>qA�<`SwpN@M_O]n����CFd XF�0GR�0��M��NFLI���/@U�IRE�84�"� SgWIT=$/0_Nc`]S�"CF_�G�� �A0WARNaMlp�d�`LI��J`NST� CORz-�bFLTR�/TRAT T�`� $ACC�aG�� |L�r$ORI��.&ǧRT�`_SF\gPCHGV0I�Ed�T��DA�Iu�5T���HK�� � �#4aԂN�HDR�B�2�B�J; �C���3��4���5��6��7��8��� 4�z�l@�2� @� TRQ��$�f��ʀ���_Uؖ����`COc <� ������3�2^��LLECA�!�MULTIV4�"��A
2FS٠ILD�8�
1��n@T_%b � 4� STY 2�b(�=4�)2(�P��9Ӱ�� 
7 $��"p��*�=`�L* P�TO���E��EXT���ы��B�ю�22�08��@��%b.'�B s�;�E� �"�E�/%ua��L��3s�08�I� Gғ�/A��⋒M�� � 87ՋC�! L�0U��� LׯpA²$J�OB6���������IGC�" dǀ���� �L�-'l��;�Ƨ4�s_M��b# tǀ�F� �CNG�AiBA� Ñ�����/1��@���0����R0��P#pX��}��$��p���t6q:Q�
2JQ�_)RB�qCTJT�Y*tJ3�D/5C�	��ǧ��@�  AzO�'л!% \�0RO0�6� �IT}s� NOM_,pn#�c���ՠTU�@P�� � ��&P���� ǨP�	ѭ��R�Al@n �3�5���
g$TF'%#D3� �T��kpU�1'�q�%�aHr�T1�E ����ң�#Ѥ�%Ӣ�Q`YNT�"� DoBGDE�!'8�Q�PU���@hֽ��"���AX��"�uTAI&sBUFφ��3!��1( �װD&J`P�I84'aP�'M��(M�)6 �&F�'S�IMQS�@NKEE3PAT�nЍp,"�"�!_MC��1)G�$��`JB����aDEC[:� [5"�����* �I�CH�NS_EMP��#$G��7�_��c�/�1_FP�TC�6S���5�`��4�q y�V�x�Kx��JR����SEGF�RAe�OUaPT�_LIN�?CPVAF�A���`�7$+�� �c_BNu�DBnrB(	,` +�Ȧ9� �A�0��AX0c`5r�D8���IX1SIZ\����D�FT�C�Z%Y�ARSa��CD@�I W\%@WX�00@L�����0�VCRCӥ�sCCw��U%@�X�1խ�2�Mdq�U�1T�XxQ"�UDѤ̣�YCk�p����4?`рf��FhE�VFf�F\a_�5F�0N�ftPX1�h���)�^Cq�+�V'SCAO��A�f�2(�(��-հ	��{�MARG���U�F�4@���1DWQ�r�0LEW�!��R�P0��o�l�"R��.� ���ϻ����%Ρ�R� HANC��$LG)��a�ǐ��̀�:��AY���u0R Mr�3�s����s4 �x3RA���sAZ�0E�tB`�O��FCT�gp�FԠ�R�0D0V ADI��O����� ������)�)�����SO�[���BMP�IDPY �1��AEQS7P^c��W��N �S!�qI��/ � �PI,?��40���b@_C�$m�K?  ?�CU0ϑuU��1�TITq�0�V�%97A."Z_\`G2 ��� �!��vNO_HEADE��!~�w�l�0��z�S+�q�R9����43 T��b�5CIRTR�0�W�X�LMt dC�gRJ�����!ERRL�X� �4�Q͠ORB$ᢳ���{�$R�UN_O�p�P$SYSР4�͠���U�EV�W�ǡP�XWOyP �5$��$SKc�"אȠT��pTRL��6̐p�P�����INDI �DJ�d�_�`�!X������PL�AS2SWAzⰰE��D!Ľ�!R\��UM�MY9��1� M|�DBO���7E���!PR~Q 
?��D��-���8 lК$f�$Q/�L�9+�����P �:Q�ãPCr��;pς�ENE70�Tq<��c���R�ECORj�=H� aO�@8$L��9$Þ"9���0F@t�JA �_Dʁ� gROS���"SK� ��rj�ׂ� 1��C��PA��>JBETU�RNA��SMR�U����CR�EWMz8B
0GNALJ ��"$LA� ���:$P�P;$P�j�{�<��!�PC���PDOR@�Q�����R�GO_AW�"�MO���p �a��DCSSp�STCY��>����0s�<�SID���2?�2M�N��OB�>&�j`I�� ? P �$@�RB�Bt�PI�M�PO��I_BY� ����TJR&�HN{DGj�@ H�`��1���0{�DSBL =��s�N�0q�W�(�LS��A��0� ,�3FB[��FE�@��N�&�)0B? �$DO�1�C�pMC��0��I�4���RH⇀W/ ?(ELE��u
r\�Ǡ(����C�q�$^�q�INK�)[�UV�L��H1A]�QoP$|#oPq#��� D �i��MDL 2C Α5��C���JoR�oR���	��g��	x��:�B�SLAVrElBING ��#��&�C�FP�@P`�p ��q�������ouСO!b���!��ID��ȃ���W��NT�V�#�VE�$СS�KI��`A�C/3	'2�IB�1J�f�1���4SsAFJ�C'_SV*��EXCLUs���NLrONL�0k#Y��x�s����HI_Vɀ^�RPPLY��R7s�H� ~�#_M�b>��VRFY_���"=Mas$IOj0��D�&��1IB�$##O��F�%LSR���4ǱI2N�.@a�P-�i$,��&AH CNf@��a5N�F3t��GCH	D�s�_�L�E *�CP��4TǱ�!�_X� G��H�TqAn���!� e�NOC
tHlB�pTQоA ~7D�$�I D $���6�-:C!$qPCF_\ NLHLC#�*�E�@K2�J��q��0x$(B� I �2_SG�` K; �ΐCUR~Л� ����A#�fЈ�(��H|(��FANNUN��@j5�CN��@�����Ѐ�YQ��$Z@V��EuFРI��L @�`�FR��	$TOT �Ч��03�ձ(5��ǠEM+�NIK�M�6�R��RA��TD{AY�LOAD���䴧R�5���EF_F_AXIJ�N���ڱ�O`=À�_
��QqO2@�`�6`
BcE�Kce� �Nh Qw1a���A8$p&aqP 09Q�a`n� �a�ӯvDU��گu�^�CA �QjR���n ,�IDLE_PWGs�e�-�V��V_�`� ����DIAG_�Rߜ 1$V��SEs�T}�6q� <zDǰR���QV�7�@SWsq�� Cp�`�1e� O1a3OHGe�aPP�IR��B>��b� ᑠ�:P�r6��x� R��u���e� Qh 6`�,�:uRQDW�uM	SG�6�A��uarLIFE��BSQ@��"Ns�=r|�Qq�=r�C8�SC�@@�Nr�YՐ�FLA�3QOV Ј�퐰��SUPPOn���"��_��E��_XP*����Z�W�� ��q�	��XZ�_A�Y2o�C"F�T(�)�;uN�9u�Q� �vn@��I{CTlS `��CACHC��ؒ`��Et#��y�SUFFI����=���b�6��	`DMS�WɕT 8(PKE�YIMAGf�TM ���SU��BQ�Jg��OCVIE}p��U; hBGL�P��?�t@W��0ʔV�2@��ST ! ��YpŤհŤ�PŤ`ŠEMAI� =��Q�%��1FAULK�WX��<�u�AX�U�Lx�pTB>PnXC�R����X��&�0���_LDEBU ����%�T���aY< �$y���S�`�`IT��BUFꗤ�r��N�!wpSUB�����C�#�z��q�SAV𵲲7p��Yчp�  VP������~t��_��ֵ�PL�OT(0���cP� M�vČ�2s�AX�S]P� Xإ�M#$�_Gs�
G��DYN_�q�PZ� <@`D���+���rM�bT80F�g�%�0DI�2EGDT_{���Q[E� GƱxQ&�C������a��ҷQ\� ��� %�T�C_R��IK�rb��B_�=�RM�^��B�DSPde�B�P� ��IM� ���ѥ5B�*pUy�ހ4g�`�M�IP�B��q����TH��y��2`T�q��HS�~�GBSC����`V��P�J��R�_D4CONVW!G4R䍐$�֥�Fsq"d~�������qSCr�T�M�ER�$B�FBCM�P�#A�ET m]C�FU��DU��b/�o e�]2CD����g�����NOa1�Q^2B;��U;��U)P�1=�C@J��1�p�u�8�z��P_H *J�L��0�� ��>P��#���1���Q����Q��a��-���7
��8��9��s�����U1��1��1��1��U1
1
1
1,
�2:
2����2��2���2��2
2
2�
2,
3:
3��3T����3��3��3
U3
3
3,
4:N��EXT-q�Q`�� �����������'_���0FDRtaT��VC0n�v�D!\J�v�REMUpF��N��OVMu�j%As)oTROVs)DT��6�*MX�,INs)����*qIND� ��
�(	�v���G���s� ȳ�|�bqDFf� RI�V�0����GEAR�u�IOYuKc"��N ��Q8aW�S�q����Z_MCMg�v�1 r߀U@��b ,H�ȱ? �A��\�0rq?�1E9p�1�����9"�c`!�P��)pR�I�5�ETUP?2_ d �P��#TDDЪa��T�@�1pGE����BAC��Ge T����(�)"��%nS�����IFI��q����@oEPT|rt��FLUI4��f �j�_�{�UR �q۱�����Jਰ1s�V`IW$$�BS�@k?x�@J%�CO?��b�VRT�yPx$�SHOUaJP�AS�SZ�m����$BG_`MQnMQ��MQ��<MQ��FORC�3�C�DATA�ag�F%U�11�S2:Ҕ1��A���ah |� N;AV}���@R��_ S���$VgISI0�SC}ģSE�07P�eV`O�a$a�B�B�A�`^f$PO�PI�q�FMR26%i C"S��b D!6�^fH'O?a?s?�&(I�:uc"_:>FpGIT_�A�TpM6|-??=DGCLF�u�DGDY'xj���DCG5��?|��1M3��jy��i T��FSJ���k P���r6�v�$EX_�q�x�q1���࿂j�p3�{5�v�Gf��6%l �� ��SWٵONA�k�QTl�h%�GR&@f�U��BKmU��O1�  �P�7`�`K�7���
�7�M�6PLOO��y�SM��`E���A� p_E m ��-!�P/TERM��n��Aa'ORIѠ�o���1GSM_#в���p���nq�P�q���qUP>��r� -�!r�m�@��)�n`G\.�@pELTX����FIo��њ0���Ʉ%�o$UFR)�$>�X����f�`OT����TA,��W`��NST�PA�T!��PTHJ�L��E��'��X�ART�b�Yp�����REL���SHF�T��ȑ��_"PR(���� �$��X��q�aE P�Ӵ�SH�I'��dU�� O�AYLO���a���@�0�-Rȑ�QR��ERV ���BC������``�@�n�@RC�1R�ASYM��R��#WJk��� E�3���B�UB������Yp��P�Ӱ���r�+OR�M[c�q��Jds�R7�p�ǐ���a����HAPTI6V�t�2MA8��������A!��A⬁H9O6Pvtu Ԯ��E,6`[`OCQ�U��1$OP!dFѩ�F9S_!$PP_ 2T�R���OUL�ȓe�@Rƕ��o���[De$PWR 0IM��ĢR_J���P�ۓX�UD�2�0��x� v@$HzhE!�ADDR&H��Gʒ-�"��6�RbMaw H�S ��	a`Z�nZ���Z����SE�ac�HSv�MN�Bx``B�F"��(�$�OL��` }�%���RO�P<a��AND_C��=�x¡�Ć�ROUP��BԲ_�0�RU�ձ1� xb0��:�`:�h!;�@��:���:�yPxbA`<B2��AVED5���E���Jcy $�P��_D�X�-R�үPRM_�RܲT�TP_=�HMaz (H�OBJ`�[D$&LE������>N`{ � ��@J�_�!T��N�S԰܄��HKRL��HIT糫�NP��al�N��%R�F)Sl��Gm�SS�� $JQUERY�_FLA��"�_W�EBSOCb�HQW&^�Ma|U�w��INCPU���QO c�P�& p�%~��%��IOLN.KB} 8�RI@, �$SL\b$I�NPUT_��$p��t�>a TP SSL��Ma~[ q����~���IO^��F_AS�rQ@�$Lf@"�fAH� a��o��@a�j���HY'+�A� U;OP�u� `� I�&�"� "s��P ����i�"��ܱ�IP_MEa�A� X� IP"����C_N
��r���qI�0s�)!��SP[B��~PBPBG�B� �@��αA� l�p{�TA��)�A6P㰔n���ؚ`U%�PST&BU�`ID�p��6P|%z�`{%�1#"w"����"5*h$I$| N�(�`��%�IRCA_C}N�  � �@�m� CY��EA 
1a<g��'7�C��x=�~#x�DAY_� (NTVA�E� k7p��w#k7SCA��Fk7CLq�!-Q��"`�A��/�$��%�5N_T�C�B� �"Y1�@���P`�A���� {!��_8�Q 2�� �$!iA�A��� $RF�R LA�B��pA�`vGUNIr�dC̀ITYb�$!&�"R��
P�s�v�CUI�URL�P7�$A��EN?�ۡ��Q����T��T_UNA2 �J �Q���$R"�J�@ R�a$P�`A��.QJ���9RFL�pA0x`
|MS5s
�UJRIe� �� F�pq�P�yRD�3$J7,��RJ8�Y7�p^2$�R�W7uF�P8�Y�QoAPHIBpQ�Sz�WD�pJ7J8ڢ�`L_KE�@ o �KG LM�!� � <�0XR��  3WATCH�_VA�Ѱ��A�F'IEL��y�0(b&�u� �`��V��V���aCT�@�f����{LDM� x4�&�_M��ΡD�1Q��LNTK����COIO���fNF��fTa�`����JvP�(������LG�d��� !�)LG_SI1ZH�9�[uMRYw� ZvFDexIYxpxl� gv|x��ZvWpf�`s�v op�v� �v�p�v���v��n�P�_��_CMD��#�Lg+�'�F$��1�K�Wp��(Vqc�bqp�opp�� p��p|�Io����pp��p�p�WpRSK`א  �(2�LN�Q���ZU��DE6�E�@`��A����԰L�n��DAU"�EA��0G 6�8�.�GH7�dQ�� BOOO��g� C
�IT��l�/RE* ��S#CRX��D����>"�MARGI��Ѐ����U�ᒍ��S�.��W�����J{GM�MNCH��&�FNb�K@��@�>�UFL���L�FW�DL�HL��STP�L�VL��@L�s�L�RES��H��h��C��@��A������U��`�򗈃��`S�G0�	�POW��������,�6�!N�EX�TUI>�I�pC0�q@.�ֳ�ֳ<��A�� o���������N�����ANA�+tAVA�I�P�Ա3�eDCS�\0b�R�p�R�OX�O"d�SA3��o�S{�֘IGNpp�0�s=��`�*A[�DEV��LLF�aZ��#Cp��`�!Tr�$fw�H� 4�b��A� �B���0b  ���+S1J�2J�3J�9r8��S�Cp� �@�p)t}��~|%�����r����Q��ST[R�9�Yr�� �$E��C�ۘP����p	�炈�Bq� L  �p.���e������j�)՟�_ � �������3������MC��� =�� CLDP[�eTRQLI�AV����FL!��lQ��11Dwa����LD������ORGQ���?RESERV(M��4M�? ��lS�� ��`�������S�V����TR	1��>��RCLMC��M��_���J ��MDB�G�Q�5`1sM�A�dU0FC�U�T�8�r%E�P�s�F�RQL� � �KyHRS_RU��b�DA0$�FgREQ6�u�$�YwOVERj �s�t��~VPU�EFI� #%G�D3uYz�ǚ \P��T$9U��B?�`�1PSI�9P	��`���D"��U� %?�( 	�aMISC�kU� d����RQB7R	 pU07P�鱎AX�b#`��EXCES�B�!d)M)@oQ��`u�d��eSC�� � HA�_I@>0P+��s�K�D���d%B_�`FLI�CB�B��QUIRE �pu+O�+2vWuLd�M�E� ��{�� �b�c��ND�g0pP����Lx� 3D;�
�INAU�T��
�&p�P8��N�r�q��!��!PS�TLoQ� 4�0L�OC��RI�@��EX�6ANG*r.a�ODA]�qrBzPbMF�b�u����c⽰m��5�$S�UPi��FX1PI�GG� � � �`c��q��c�
�c�@ ���5I��EH��TF5 0t�0�TIl`C����pM!P� tV�0MD�AIB�)�FX��D���GH�0�Q�DGDIA�Q�C4PW�P�D0ѧ��ED@�)qOjS��pP� �CUppV	P��.W�Oؑ_ � �`{Еӿ3 4r��pB|XP|^r����PP{X�KE�T`e�-$B8W�oV��ND2��Pc��Q2_TXl�XT�RAX��R���� L�O:���d"�g�CR.f&c�2R�R2h�� -�a�A�� d$OCALI��uGF�:jg2F�RINb�ncw<$Rx`SW0��ܨc��ABC�8D_�J�P{!.�A_J3:�f
�b1SP� P.P�d�m3�mHQ9�
.#uJ��3un���O��IM���CS�KP��bt7�?�btJA���Qb|�uyu�u�w��0_AZ��/q�qE�L��.r��OCMP0�3���RTE�s� e1�0pe�1����� �Z�SMG�ՠ�@��JG��SCyL��5SPH_��� ��f���.u`R'TER�`nc�k`)_E���b Aؐ��̯�DI�qQ�23=UdrDF  � ŀ�LWʈVEL��IqNx���_BLX�.��Yq/J��������IN���]`��CR9�ْ.�8�6�_T �F�a���W �^�"�k���"�DH���P\a���$V0w`3_���$=���~&�$��]0R�6S]`�H �$�BEL�pm��_A7CCE�� 	����IRC_��q�@�NT��$P)S���LЀ�0M� ��9�.��1G�/��Q����$���3S�T@�_�G�ؒ�����8�_MG}DDء��~FW��@���$����DE�PPABmN[�ROg�EEˢ K�B����qK� �~Ѐ$USE_v`��P$ CTR�Yh4�ꐪ� ��YNgAA鰢�Rp�A��M:�NQ=�ҠO�v�ϴINC(T�1�����\Yq�ENC��L�A`.K���H�IN��aIS�8ť@O�NT�>�NT23_Ȃ~�f�LOـ~|�� I � #��΀#$ ��h���#"CQ�M�MOS�Iݡ<"[P�����P?ERCH  �ó�� �Ǚ1��lA�­�lA�w�r������PsAS�E�L��Ps7'OwN�p@�ʄ֟�TRK��R�AY"c?�!��S���ոӔ0�v!��P MOM鲎"C�HP$��jg�ӆ�g�T`D�UXp��S_BCKLSH_CS�F�:  �ƴ ��-e��o깱>�uCLALMJ�@8�Њ���CHKep�@>�TGLRTYp@�S�8ėE5�A_�3��_UM3��C3�Z��� LMT�`_L G��s%��A0�E*�K� =�)�@�F�@�p9N�L��)�PC��)�H@8� ܥ��CMC�U�.�CN_�bN�S��&;sSF���V���A�.ǃ���S�/��CAT��SH�3�b� � ��/�/�eT�i�٠3PA���_P����_fpZ�����eq������JG�0��ӀO�G����TORQU ~��e���� �e"�� �B_W���ّ�aʓ`Г`IhI
vIГF�0S:r�,Iq�VC�0!%��1�ڠ��q�J�RK�!"&<PDB�X�MtS<PM0_D9Lʑ_�GRVg`$0ʓ`$ГA!H_%c?#���*COS�+�p�(LN# �+��$ʐ�)�=��)��*�,�<%Z� ��A!MY�!:8�"��Q�+[9THET0��NK23Г�2ē�� CB�6CBēCz`AS�A�2��1ʓ��1�6SBʓ�2�5GTSkqZ�C�a���&�J�#$DU���h�6Bjb��EG�Q�%�_��xNEht�s�K�������y1A�}5�E�G�%�(�!LP!H�%�B^ńBS��C �%�C�%�B6!SZ(6��@V�HV�H���LV��JV�KV
[V[V*&[V4[VBYH�H�F��R�Md�X�KH
[H�[H&[H4[HBYOJ�LO�HOsi�NO�JUO�KO
[O[O&[O4[O(6F�B�1y��%t�GSPBAL�ANCE_J16sLmE�0H_}5SP>���&^r�&^r�&PFULCbx�rqw�r�%K�{1��UTO_�����T1T2�y
�2N���V��tM��ыpPi@Z��	�Tu�O��|�QINSEG����REV���G�D3IF��p�1�U���1�y OBK���j#��2,V���I$LC�HWAR4���AB���$MECH`�1J0��ǁ��AX���Po����G���p� �
�?�0�ROB���CRS�#���	 � �C�_�T �� x $W�EIGH��w $ȹC\�� I����IF�v��LAG����S���:���BIL��O1D�Ы�s�ST�s�P:���t��N C�
L��P�
������  2���x�DEKBU��L|�Ē5@OMMY9C�9�N��$�w $D|� ��$�� l1 _ �DO_:�AK�� <_�ޖ�p�ᰱ��@B����NJÁ�_ԍ��� ˒O�� _�� %�T7��?��TL��F�TI�CK����T1N�%֣=�ߠN���pu���R\ఱ��񥩂��U�_PROMP��E�B? $IR"��p��8�X�w�MAIF h���Q�_��O��X���°RU COD��FU����ID_�����8�2�>pG_SwUFF� ��4��X��DO��/�������GR����Ѵ �ݴ��赩���-Ѵ�U�퐱_�H�_F�I�9G�ORDf�� R��36s��H®�N�$ZDTΚ���ˑX���4 *W�L_NA���ߠ���DEF_I�ȡ��������������������IS�m@# m�|@�0������6�4���DP�p?�f��DO@p>l�LOCKE�˳����2�Ѳ˰UM е��Ѵ��Ѵ��Ѵ>� ݲ��ܵ��ݴ�ݲ�� 2�2�賴��赡��@���9�w�͸��P}�  Դ�,т@F�W�ر嚨���TE��Y��� ��LOM�B_����0s�VI]S� ITYs�A�}O��A_FRI�s��~�SI,��naR�ܠ7��7�3��s�WB�W�Q �% _���EAS{����P| x�W�8�45�55��6|�ORMULA�_I��G�ǵ� h 
�7�C?OEFF_Oá&�H)á�0Go{�S���5�CA�p:�L�ˑG�Rm@ � � �$���rv�X��TM�ד��ɢ�ӭ��ERI�T�Ԑ�퐳�  �rLL�p�SΛA_SVk��$���퐴.0��퐵 ��SETU,�MEAG����t�ˑH�>L�� � (� ���lقl��Dw��ߠ�ќ�}Ԃ]d�����y��G�xг[@��k�R�EC[�q��SKy_Apy� P_�?1_USER�q�2�$��*4 �qVEL@� ��-"!%��Iz���p�MT��CFG>��  �]�=OςNOREJ���~l"�OPWOR�@� �,B�SY�SBU�P�SOP(�!��T�*U�+X�1P��K"�%PA qX�#˂�OP�U����!}����� IM�AGz�� d�IM� 5IN���"3?RGOVRDfP�#	 �!P� 3 �|@g�hl�i5ЂL��BT:B>lPMC_E���!��N�`M�2��1��>�H1SL|p��{ �R�OVSL�S��DEX\���5a@��8_H0�7�I0��3��3GH�4CC�����5CAGI0_Z�ERl!�2:��O @ _C�O��RI����
�Fg��I��A�A  �Z�EGA�� H_�̀Ð�ATUSk,�C_-T31DX�FB� �F��ApV���C���� Dc�� �2�B�P-�`�AM�- �r1XE�@ x9RMRTvC�}@`���@UP�H�&�PX�;�V�1�3�7R��PGY%�� $SUB�A�E��A�CJMPWAIT�P\C�ULOWςFʡyM��ЁRCVF_�X�ς�QRE`F0���CF@RLς�<gIGNR_PL�C/DBTBÐP*�Ё#BW�2dt U��1e�IG�!!��qҀTN�LN0f�bRT{3N�O�N!��3PEE�D�P�3HADOWxÐ΃t ERVE�3��d�2�Q��SP�p � L_�瀼��`1�tUNq��[p�QRTPNCLYw���A��1PH_PKT�Z#�b"RETR#IE�Cx"�"P!WpvD�FI_r� �R��Zp�t 2�d D�BGLV@cLOG�SIZ܁�ZpaU�m��tD�c�`_TX�τM��C�B�EM��}R�s��ˆCHEsCK~`��PL ��� 0@vx9�A3LE�Qx�PA�Ў�����rIP�b��
AR�r��N�=��b�@O��b��AT�� xc��v�pل��1scUX� ZBjQPL���Z$� $d!��SW�ITCH�rE�WO���A�R�LLB���� $B�A�DvӞBAM��@.�C=��A,�J�5�`N!Y�6_��_�KNOWO�u�L0UF�AD/�c 
pD ~��PAYLOAq�9ී_�A���!��Zʽ�L�Aj��LC{L_�  !4���S�?!�]2�F��C� ��p�� I���R� ��W�@P�Ḅ�� _J�b~�_J��� !SPTAND�q�������~!��P�L�AL_ Ȕ�
pA�B�1��C�D��E��J3ܱ�Ŧ� T PDcCK�0)ҞCOMfH�PHգ�BE.��կ��X|a�0� � ��`��D�_1��2�DMA�R@Q��������:PR�TIA4ù5ù6�MOM��ϳ�ܳh��V B`ADϳp�ܳ��PUB�0R��@�ܳ@�:�+������ L$PI�4�at�!��=ATܙ��I��I��I�À����\��ơQ�ƬQ$RO�c��E�cHIG��ce�d4� �de9`.`4�j�C�9axR�9aeSAMPHP�=���4ק�eN��� &��� ��!"�Ԁ�P���`���ٔ�!"R���ȴ�Տ�m���IN 5����<�X�3�b>��~�U�~��GAMM�*�S�A���qGET�!�FIO��c�>"
&WIBF�bIl�d�O$HI���A�@$!"�E;� �A�=�.�LW�[�R�=���.�X֚`ǡCheC�HKV0�@�
�I_�Й�>"1�r�v�$������1���ţ ��$�� 1����IRCH_�D#��P$d�LE@;!!�At^�< ʧ`_MSWFL3dM��7SCR�X752�p ��O����F�ϰ�ٰ�	�`��SV#��;P�pCUR�#f�pSAA�n4A�NOb�C�A�c�A ��r�ȟڟ�Ȯ�����������DO�aA ���q���
�.ؚ">��^�j�?';%��� ���l�Mq�� 7� ��YL��r�$����p�%�r�'@`�@	�"�#r�(0� �@a7QM_Wp�" �"`��#��s!MG`�+��'ġd�4���5�Rl�M2wB� �8�q� �4$WQ0�5ANGLa�Q0:� O2A�O2H�O2�X`;�ANo������sw�XGp	OI�v�Z�5l�`rķ� ���OM ������ư�p�g^�LNKl�b�_�R� |�HN� �Fܳ�F:�NȺ�G�F�����i�o"B�O  �DP����PMON_QU��� � 8:�Q�COU:�QTH�|`HO�"FPHYSf��EST�FPUE1Pt7�PO�T�  gp�P`�bRUN_+TO�#UpO!��� P���U!e#I�NDE�sc�GRA�� ܀� 2� NE_3NO�T�UITj �Q^sPINFO�erh�[a�"��1OIb�� (��SLEQ@%�.a�.`�VrQS���p�� 4:�EN�AB}2�PPTIO�N���d�g�dbcG�CF�q� @:�JX0v�R���R�h�hq�o�dn"��EDI�T� ��p�0K�E�&�$�E,�NU�wxAUT]uCOPYE�!�6|�i�M�N@pD{��PR�UTq2 GrN�`OU �$G�R�t'R_RGADJq�y�X_� I\�0�v�0
�vW�xP�x� �v=���pBbN��_CYCz}2i�RGNSge9� w�LGO����NYQ_FREQ�W�W���\����SL�򐞂T��q곉�&�CcRE��QS��IF����SNA��%��_}GjSTATU�@<j�WMAIL�Ҁ�yIuATLAST偼�.�ELEMka�� ���vgFEASIxa?"��� � �&� JE��b!���I�P���S��IQPyz�AB$�a�E�PA�V���~�����X�U_�!�V���ǖRMS_TRt�v�g ��3^�Bb �Ɣ �00��3�݊@	Q� 2� d�4R�7��� 6��.0 �!��b���NnDOU�SbN�c�0�PRd l`�5bG�RID�Q�cBAR�S%�TYyc�rOT�O
�q� �Q_"��!�pݢ��O�0hd�� � � �@P�OR�S����SReV��)&��DI_T��?�R��\��\�Q4Z�� \�6Z�7Z�I8>�(QF��ka�~P?$VALU��4�7�5�qQF4���C !teX�Q����1�`AN3�́R�pa�5�TOTALX�Ӱ1A�PWI�I��>W�REGENU�j��CXӘ�Sa�Q�,PcTR��W�U�_S7��j��cV�q�d�¢b��E샩�KQ4��R,pn�V_HƠDA,C���S_Ye�2m��S� AR,@2� }�rIG_SE��������_�P��C_�Ѧ$CMPp7��D�EtKБ�I��Z���\�Ba��ENHA{NC2Q� p$��ve̂ ��INT�=�g�0F�S�1MAsSKȃĐOVRQSP#P��H@��vầ�V�e ���pb��V���>Ѧ�PSLGT�ka�`=n��02?��H�S�"����U��2��TE�0İ�#���o��Jb�]}�IL_M|��w���@TQ,P��Q͐ԑ�"V2�C@�P_h�VJ�Ma�V1`��V1n�2}�2n�3*}�3n�4}�4n�#���!"#�`���!"IN	VIB<0:�' T!.2*263*364*46p:����Np�T �$MC_FOPd�$ LBN��5�MbnI�Ӳ~� �@�5B��� KEEP__HNADD�!�$���	C�1��ݡ���O%Q�zp�p2 ��REM%�G� �JafU���eHPWD w �SBM�~��COLLAB.4����3���`IT�3��0&rNO5AFC�ALt2��4� ,�7`FLz0��$SSYN� ,M�@Co���V�UP_DLYzq�~RDELA= �H�ɂYPAD,A�:�QSKIPS5�� ���PO�0NT�!g P_�P�R�' �P�2g��'���)�a�) s��*���*���*���*Ч��*���*9�q�RAhd� XJ�'����MB3NFLIC��S[0T�US����WN�O_H[ DHq�2IuT�r<0_PA�P�G�� ����U�ҐW�`�6M���NGRLT= �Q�q����p�����1�T_J�!�6BbAP��WEI{GH�SJ4CHxP��4OR��4$�OO+���d��6J	���aAaA��nCIHOB`�L`���J2s0q�pcX��TV��A�Q5��A�p��A�Q�  ��RDC��� ��
pR�cR0P9�"R����JIR�B9�RGEp�`c��C��FLG7p�PH�d9�SPC�S��UM_�@��2T�H2N��_@�A ?1� �s0ݡ>4� � D����\I��2_Pd2�S�S����]�L10_�C{��1�T�� ��p$�P2�Y��C �;�� a�D��aZ��Q�C7c���h���`�U�МP� }P��DESIG�R.V�VL1�Y1�VTcvg10a_DS��l�92EFOp11q� l� ��!��ATC�t��_��bIND����aOp9�x�b�2HOMErS �Q�a2�b��o��o�o	-a �d3�b�Pbt���S aa�a4�b�������'�?p�$�$Ch�SBP��i�ā77 ���	�SI"��π�Z�$AA�VM_WRK 2� ą �0  �5�ˁ�%��H� H�	k�\��7ŀ!�m�������[�Ν�ڟj����'�/��B�S�`�A 1��? <�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D� V�h�zߌߞ߰����� ����
��.�@�R�d��v��?�C( AXL�MTBP���X�  d��IN����WPREoPE�������_C_��O  ��� c��� �I�D ?ą�� 8�d�^�p����� ����������9�-a�0��J��UPb���4  �IO�CNV_lP�� ���P}�0��T�>�V@�  1 �P $��畑���ŀ?�L�� $6H Zl~����� ��/ /2/D/V/h/ z/�/�/�/�/�/�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFoXo jo|o�o�o�o�o�o�o �o0BTfx �������� �,�>�P�b�t����� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�D�V�h� z�������¿Կ潝��LARMRECOV M�����LMDG -�� L>�_IF� ���dF�ILE-066 �UD1 Ins General���isk 234 �1 mode J�1 at EOA�T chg,G1,A1) 11���  uted VPL���������!��3�W�, 
< �BA���8 �ߍ�A�UTO�� WORCLDo������ R&�UPPROGRA�M LLET_R�IGH����ABO�RTE��QNGT�OL  �	 �A �Z�h��P�PINFO H� Gƞ������}�  T����-� ��-��Q�;�M���q�`�����������+� 1CUgy�������3�PP�LICATION� ?������Han�dlingToo�l�� 
V9.?10P/23z���
166775�57H745891��G264H=>O7DF1C�ޤ�None��FRA� 0���_ACTIV�E�  R�  �#��MOD �]�P�%CHGAP�ONL?/c�V OU�PL�1p�� �� �/�/�/
+CU�REQ 1	p� U ��,�,	? $594.��/??+?�=?O?a?�?�?.�;�"�%�4��"�:HTTHKY�?�?�?�?�? 4OFOXOjO|O�O�O�O _�O�O�O__0_B_ T_f_x_�_�_�_o�_ �_�_oo,o>oPobo to�o�o�o�o�o�o (:L^p� �� ������ $�6�H�Z�l�~����� ��Ə؏��� �2� D�V�h�z������� ԟ��
��.�@�R� d�v���������Я�  ���*�<�N�`�r� ����𿺿̿޿��� �&�8�J�\�nπϒ� �϶�����������%�TOC�/1#DO_CLEAN`/$���NM  H� �/����	��-��.DSPDRYR��&%HI= ��@�ߙ� �����������)��;�M�_�q�(MAX@~�7��o'��X~����"�"PLUG�G~ ׋#/%PRC*P�B������z����O��Y�k�SEGFW K5GR���߀�����LLAPv��35GY k}��������/R#TOTAL�����R#USENU
v �+ d�h/�� �RGDISPMM�CU ��C]��@I@k�$Ot���a�#_STRING� 1
O+
�kMH S*
�!�_ITEM1�&  n-
??.?@?R? d?v?�?�?�?�?�?�?��?OO*O<ONO`O�I/O SIG�NAL�%Tr�yout Mod�e�%Inp�@S�imulated��!Out�L�OVERRs� =� 100�"In� cycl�E�!�Prog Abo�r�C�!�DSta�tus�#	Hea�rtbeat�'MH Faul0W9SAlerCYsOa_ s_�_�_�_�_�_�_�_o z��+z��/ oTofoxo�o�o�o�o �o�o�o,>P�bt��oWOR U �+�qDo��
�� .�@�R�d�v������� ��Џ����*�<�N�PO�+$Qt��{ ]�������͟ߟ�� �'�9�K�]�o����������ɯۯ�o�DEVw�����?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ�>��PALT0m�� ���������,�>� P�b�t߆ߘߪ߼����������(��GRI���+`���:��� �����������*� <�N�`�r�����������N�F R0mx��� ,>Pbt��� ����(:�L^p��PREG �Ω����/ /*/</N/`/r/�/�/ �/�/�/�/�/??vM��$ARG_�pD ?	���W1��  �	$vF	[�k8]k7�vG�9J0S�BN_CONFIQG�@W;�A�B�1��1CII_SAVE  vD�1�3J0�TCELLSET�UP W:%  OME_IOvM�vL%MOV_H8@$O*OREPuO�@:UTOBACK��1W9�2FRwA:\� �O,��0'`P��H�� �K�0 �18/07/�10 22:%P18��8�6_H_u_l_�L���_�_�_�_�_oo���_DoVo hozo�o�o)o�o�o�o �o
.�oRdv ���7����p�*�<� �  �A�_�C_\ATBC�KCTL.TMP DATE.D�����������ˏ�CIN�I���E�6�CMESSAG�0��1_0��3�1��ODE_D�@�6�$�O�,�ޒCPAUS�� !��W; , 	���0�� ���k��
�����!���x|����(�,		 ��W5��Ɨ���П� ���@�*�d�N�`��������̩_�i�TSK  o��A�1��J�UPDT#��d�9�Z�XWZD_E�NB脸:B�STAp�W19�I1XIS�0?UNT 2W5�1��0� 	 �={�����pP����}��eӖ��� 
Z	 x�� L�  #�� .5 3�q����	�̱�h�� <�+=� "U&R'�Ϳ���
�4�p���}π�MET �2��3 P��H��HY�|H�9{E�#UH?S�AH�%;���@�|C?Nl��?�<�TN�>���?������SCRDCFG� 1W5�A ��5�2m�A�S�@e�w߉ߛ��O�U�9 .������!�3�E�� i��ߍ���������0N��B7�AGR��-�XM�&�^�NA>@V;s	�D#�_ED��1��I��%=-d�EDT-�RJ���� ����B����2�_����.D ����29����<����b� &�J��3QK �`R���.������4�A/e w�e/�,I��/V	5�//�/1/w�/1? x/�/ ?�/��6i?�/ �?�/w�?�?D?V?�?z?��75O�?�O�?w�^O�OO"O�OFO��8_uN_���*_�_ �O�O�__��9�_=_oa_��_ao�_�_Po�_��CR8pO�o �o�M�o+ro�o�o�&�s�NO_DEL�2�$�GE_UNU�SE0�"�IGAL�LOW 1V��   (*S�YSTEM*��	$SERV_G�Rj���pi�REG��u$���pNU�M�8�&�PMU|�p�LAY����PMPA�L6�CYC1�0r~��o�s���ULS��l����i��s�L����BOXO{RI�CUR_�~&�PMCNVa���10��M�T�4DLIM����	*PROGRA�tPG_MIs������AL}������Bڟ�~$FLUI_RESU��(����C|C`� r���������̯ޯ� ��&�8�J�\�n��� ������ȿڿ���� "�4�F�X�j�|ώϠ��x&�LAL_OU�T �{E�W?D_ABOR�����ITR_RTN�  ��=�
�N�ONSTOj�5�� �xCE_RIA3_I�p5�~�A��h�FCFG �V�~�u���_P}A��GP 1�����������C�  >@�@�@�@ྪ@��@��@��@��z@��@��  D��+D|�|�8�S᪓�@�@��@���@��|���D� �D|� ���pD3���=|�F��j�DYe��?��h�HE`p�ONFIU����G�_P-�1�� }uV�8�J�\�n�����������KPAU�S�1�~� ޛ� �	�����|���s�����ݍ��?b�� x��Ϻ� 0�Z@j�v ������ �DVh�M*�NFOw 1��� � 	�ߝ���������X�S���ؾ��¤@h����1k D�z��?�EC2���ݖ����F�B_���h�O����ߧ�!LLEC+T_��y� �9'EN}�5��U"!�NDEA#I'��s>r1234567890�'9b�qp�ҧ/�&.c
 H��.c)�/?�l�/?^? ;?M?�?q?�?�?�? �?�?�?6OOO%O~O IO[OmO�O�O�O�O_ �O�O�OV_!_3_E_�_��ͅ$�q2I+ ���X+�"IO  �)U!.g4�o.o@olRo�WTR��2!�]�(��i
{_`n���"�]�j��]&_MO�R�R#�� ?� 9B����u�y +O=s�{�b��*�Q$�m,��?����HW��q��K�ty���%P"&I/�����.�@�t�
�r�/'��
�e�i@���|��c� ��a�hPD�B�p(�̉Tcpmidbg���1�&*�:�^��p�]�,(����^����l�o���K��m��Ɵmgڟ3������f"�{�<���Pu�d1:��ɯ�j�D�EF '4c)���cّbuf.�txtԯ"�կ��_KMC�c)���Sdg�H��d*V���ԕ���/3��C� B�!��C9Ca�C�A֨l�C2�IC�2��D�n�D���MD9�CL~�	D�mES��4�F,��F�� F�iE�{��
�Gb�7�Nkr  uD��w,�\�rШ�cĽ��j�`��c�`�x��۱��Cf@�z�����^�D��E�H�D��D{��F��3ES�F��I3��F��E���E{�H��F{�G�����_  >�3��C�r���n�ѧ���5ِ�ᧁcr��A�q7�=?L��<#��ea�X߉�@�RSMO?FST %�X���P_T1w�DEw -����a,;��;�Q�s�m��?���<�M^<�TEST�+��RC"./vC���A�7������?ї�B�લ����C��������:Sd��b[�I�#/e�)?��r0�m�$r��RT_�PROG ��m�%3�S�X���PNUSER  �r%��f�KEY__TBL  �����	
�� �!"#$%&'()*+,-./�'�:;<=>?@A�BC�GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������-���͓���������������������������������耇����������������������Q'�LCKq�m�h��q�STAT�Y�_AUTO_DOo&ul��INDj$D�8!R����"-�24�!# STO��  TRL)�L�ETEo'{_S�CREEN ~�jkcsc"�UlMMENU {11� <B� A�	/X��/G/��$/ J/�/Z/l/�/�/�/�/ �/�/�/7?? ?m?D? V?�?z?�?�?�?�?�? !O�?
OWO.O@OfO�O vO�O�O�O�O_�O�O _S_*_<_�_`_r_�_ �_�_�_o�_�_=oo &osoJo\o�o�o�o�o �o�o�o'�o6o FX�|���� �#���Y�0�B��� f�x���׏���������_MANUAL\p�ZCD��2�ِ���R��gߗ�?G|(�g�L�@�3F�G B��7�z��7�~0��$DBCO�RIG��	�_E7RRL/�4V��a��>�P�b� 둟NUMLI*�W�g�m�
�PXWO_RK 15V�-��¯ԯ���
�[�DBwTB_� 6�ԕ�b�t���DB__AWAY��/GCP m�= �^��_AL*��^��Y�o�m�&`�� 1}7�� , 
��M�e�(�v찅����ݾ�#�_%MI��l�@@�4��ONTIM��&m��Tƪ�
����MOTNENDu����RECORD ;1=9� �"�#�G�O�����#�m��XECUTING R�&�8�J���T�{��� ��Ը�������]�� ����H�l�~���� ���5���Y�� �2� ��V�A��������� ��k���
y�.��R dv#��? �*�N�r �����;�_ /�8/J/\/n/��/ /�/%/�/�/�/?/ 4?�/-?�/|?�?�?�? !?�?E?�?i?O0OBO TO�?xOcO�?�OO�O��O�OeO)�TOLEoRENCk�Bȴ��y�L���CSS�_CNSTCY +2>���a�_���l_z_�_�_�_�_�_ �_�_
oo.oDoRodo�vo�o�o�o�oGTDEVICE 2?W[ F�#5G Yk}����#��HSHNDGD @W[��Cz�z��JQ_LS 2A�m� G�Y�k�}���������IRPARAM �BY�k�v�5��RB�T 2D��8��<ذ C�;P��ª  �:;P�Q��@W�F��E�?�
�Q�HZ�Ԑ�M\^��@��F�x�M�C�J��8P �V�͐ŌU��;�B�8J�6UŅD�@����;���h��\�X�ńc��ņ���Z�l�~� �������د�7��� �2�ŅC�,�D�
�D0N�� 	���9M<A�+��A��,A����A��A�U2dŊ��Cs���B����4δ�Ō���|%�Bwq�B�0N�B��QB�>_C񹴿ƿؿ����? ��� gp� ~�H�ō-� O�a���I�wωϛϭ� �������B��+�=� O�a�s��ߗߩ����� ������'�t�K�]� ���7�������
��� .��R�=�v���cϑ� ������������< %7�[m�� �����8! nEW�{��� g�/�4/F/1/j/U/ �/y/�/������/� �/�/B??+?x?O?a? s?�?�?�?�?�?�?,O OO'O9OKO]O�O�O �O�O�O�O�O(_�/L_ 7_p_[_�_�_�_�_�_ �_�/�O	_6o�Oo1o CoUogo�o�o�o�o�o �o�o�o	h?Q �u������ ��R�d��_��s��� ��Џ�����*�o 3�E�r�I�[������ ���ǟٟ&����\� 3�E�W���{���گ�� ï�����X�/�A� ��	���Ŀ���ӿ� ��0��T�f�A�o��� �υϗ��ϻ������� ��b�9�Kߘ�o߁� �ߥ߷��������L� #�5�G�Y�k�}���E� ������$��H�3�l� W�����}ϫ����� �� ��	V-?Q cu����
� �);�_q ����/��*// N/9/K/�/o/�/�/�/���$DCSS_�SLAVE E�����!���*_4D  ��.3CFG �F�%3�d�MC:\� L%04d.CSV�/��{?  ��A V�3CH�0z��/�g>�?�?�  �g6��1O�9A� �J(C�;g4���0�7,4RC_O_UT G�+OB��/_C_FSI �?�) :Kg6�O�O�O�O�O __F_A_S_e_�_�_ �_�_�_�_�_�_oo +o=ofoaoso�o�o�o �o�o�o�o>9 K]������ ����#�5�^�Y� k�}�������ŏ�� ���6�1�C�U�~�y� ����Ɵ��ӟ��	� �-�V�Q�c�u����� ��������.�)� ;�M�v�q��������� ˿ݿ���%�N�I� [�mϖϑϣϵ����� ����&�!�3�E�n�i� {ߍ߶߱��������� ��F�A�S�e��� ������������� +�=�f�a�s������� ��������>9 K]������ ��#5^Y k}������ �/6/1/C/U/~/y/ �/�/�/�/�/�/?	? ?-?V?Q?c?u?�?�? �?�?�?�?�?O.O)O ;OMOvOqO�O�O�O�O �O�O___%_N_I_ [_m_�_�_�_�_�_�_ �_�_&o!o3oEonoio {o�o�o�o�o�o�o�o FASe�� �������� +�=�f�a�s������� ��͏�����>�9� K�]���������Οɟ ۟���#�5�^�Y� k�}�������ů�� ���6�1�C�U�~�y� ����ƿ��ӿ��	� �-�V�Q�c�uϞϙ� �Ͻ��������.�)� ;�M�v�q߃ߕ߾߹����������$D�CS_C_FSO ?���?�� P ��\����� ����������"�4� ]�X�j�|��������� ������50BT }x������ ,UPbt �������/ -/(/:/L/u/p/�/�/ �/�/�/�/? ??$? M?H?Z?l?�?�?�?�? �?�?�?�?%O O2ODO mOhOzO�O�O�O�O�O �O�O
__E_@_R_d_��_�_�_%�C_RPI<�N�_�_"oo �_;��_.owo�o�o(�SL�_@l`�o�c�o  $;HZl� ��������  �2�D�[�h�z����� ��ԏ���
��3� @�R�d�{�������ß П�����*�<�S� `�r���������̯� ���+�8�J�\�s� ��������ȿڿ�� �"�4�K�X�j�|ϓ� �ϲϽo�fYo�a�o�o �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg y������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/�/�/�/�XNOCO�DE H]e��GkPRE_?CHK J]k� �A � �< �� ]ee?w?]e 	 <Y?�?�?�� �?�?�?�?O+OOO aOsOMO�O�O�O�O�O �O�O_'__K_]_7_ �_�_�?{_�_�_u_�_ o�_oGo!o3o}o�o io�o�o�o�o�o�o�o 1CgyS�� �_�_����-�� �c�u�O��������� ᏻ�͏�)��M�_� 9�k���o���˟ݟ�� �����I�[�5�� ��k���ǯ������� �3�E��i�{�U�g� ��ÿ�����ӿ�/� %��e�w�ϛϭχ� ���Ͻ����+��O� a�;�mߗ�q߃����� ������!�K�A�S� ���-�������� ���5�G�!�S�}�W� i������������� 1gyS�� i����- Qc=O���� ��//�/M/_/ 9/�/�/o/�/�/��/ ??�/7?I?#?U?? Y?k?�?�?�?�?�?�? 	O3OOOiO{OUO�O �O�O�O�O�/�/_/_ �O;_e_?_Q_�_�_�_ �_�_�_�_o�_oOo ao;o�o�oqo�o�o�o �o�o9K_3 ��m����� ��5�G�!�k�}�W� �����������Տ� 1��U�g�]O����� I�ӟ埿������ Q�c�=�����s���ϯ �������;�M�'� Y���y�����˿e�׿ �ۿ�7�I�#�m�� YϋϵϏϡ������� !�3��?�i�C�Uߟ� �ߋ����ߡ����/� 	�S�e�?���u�� ���������=�O� )�;�����q������� ������9K��o �[������ �#5AkEW �������/ 'U/g//s/�/w/ �/�/�/�/	??�/'? Q?+?=?�?�?s?�?�? �?�?O�?�?;OMO'O qO�O=/kO�O�O�O�O _�O%_7__#_m__ Y_�_�_�_�_�_�_�_ !o3ooWoioCo�o�o �O�o�o�o�o�o )S-?��u� ������=�O� )�s���_������o�o �����9��%�o� ��[�������ß�ǟ ٟ#�5��Y�k�E�w� ��{���ׯ�ï�� ُ�U�g�A�����w� ��ӿ����	����?� Q�+�uχ�a�sϽ��� �������)�;�1�#� q߃�ߧ߹ߓ����� ����%�7��[�m�G� y��}��������� !���-�W�M�_ߍ��� 9����������� AS-_�cu� ����= )s�_��u�� �/�'/9//]/o/ I/[/�/�/�/�/�/�/ ?#?�/?Y?k?E?�? �?{?�?�?��?OO �?COUO/OaO�OeOwO �O�O�O�O	_�O_?_ _+_u_�_a_�_�_�_ �_�_�?�?)o;o�_Go qoKo]o�o�o�o�o�o �o�o%�o[mG ��}������!����$DCS_SGN Ke�M��w@5a�07-NOV-�20 00:43� �10-J�UL-18 22�:49g�����? Q=�����������R�S]����Zo��5�����  9�VERS�ION E��V4.2.10�ϋEFLOGIC� 1Le?�  	����`)�`8��PRO�G_ENB  ⢄ ���Y�ULSOE  >�q��_ACCLIM����s����W?RSTJNT��M�;�5�EMOb����u�
�ݐINIT �M�jזOPT_SL ?	f��
 	R5�75��C�74H�6JI�7I�5��s�1m��2I�*����&�TO�  2�����V.��DEX��dM�����PATH �AE�A\AOA{\ C�IMG\��]��$DHCP_�CLNTID ?<� � *������؂IAG_GR�P 2Re? ���`�E�  F?h� Fx E?`���D�����B�#  Ϣ����A�~/�Cf  Cyj��Y�dCj�qߪB�i����mp3m6 78�90123456����`�  �A�ffA�=q�A�  Aх�A��HAľ���������A�c�������@����g�Ap�����A���g�B4��� ��2���
����(�A�A��
=A�B����A��
A�Q��A�������� j�����j!�	n5�_�{A�Z�̶���ZѾ��������A����������h�zߌߞ߰�6�EG��A@��:�RAU5Z�/��)��#F�Z�b��������*�<�6�Pz�AJ���Y�?��9p�A�3\)A,��A&����~�������4�cF�]���AW��P��J��C���<Z�4��-Z�%G���0�B�T�6� %�
	n��?Q��% o�w��Yk� )M_�kc��Q���i������=�
==�G���>�Ĝ��7�'Ŭ�6�7����@ʏ\&��p�$%��@�Ah��/ A��<i���<xn;=R��=s��=x<��=�~Z�;���|%<'�'������?+ƨC��  <(�U��� 4"����&�C���%��\က?� �?�?6?H?h�$ T?~??�?�?�?�?�?��?)7L?S��FB$�/Eͽ,�4OG�ΐ
Ա��iD�L�x�CA��GX�j�|�챤��O�L���Oʹ�%_sN�ED  E�  �Eh� DQPXR :_���_���u�_�_�_@��q_�_m_o�K4o�:b��D�|-��0ݎC3u|����À�B�T�o�o o�o�o��o�o�o��E}��?�"� _�r>��>imߴ��Y<�=<�{Du;ě�Pu���CT_CONF_IG S׷�>��eg?�ʱ�STBF_TTS��
q��s�������v9�MAU��f�x��MSW_CFtpT�׻  ΌOCV7IEW�pU�����_Y�k�}����� ���rG�܏� ��$� 6�ŏZ�l�~������� C�؟���� �2�D� ӟh�z�������¯Q� ���
��.�@�ϯd� v���������п_��� ��*�<�N�ݿrτ�`�ϨϺ���\|RC �	V�5�r!h��^�9߀(�]�L߁�pߥ��tS�BL_FAULT� W�����GP�MSK�w��hpTB�R �X��>��q��o�F�X���TDI�A	�Yxy��s�M!UD1:� 6789012�345��rM!��P (�����	��-�?�Q� c�u�������������@���F��	�"
��<Mt�RECP���
���������  $6HZl~ ������#�52/��UMP_OPTION�p��R!�T�s��s%PM�E�uf/Y_TEM�P  È�33BȈp� �A� �$�UNI�p�u�!��Y�N_BRK Z�2��EDITOR�X!^!�/2_j EN�T 1[��&�,�&JR_SET�UPPROGRA�M H�pmpHEC����&HOME JACKPO:0�IGh?�u&M�AIN�?�? &?PICK_�?�?w#&�:LEF�p��?��&PNS0�001 OSE �E �?x8CLA�V CL<Or<&?GRIPPE�gB�nO�&X0CA�LICRA["] T��O�CCAMEA�BB�D�O�r&��H�C�@�O�p&PLACE�<$_�p�_�0=ZBHP_�pd�&X1HIP FTH�BE�A}_1W4�A�_t=ZERO �9@PALLET_�H�_z6<PSTI�C_�_�\/&C�LEAR_IO  �F�p�4t<gT dYeYo��&	MID_P�OI@0$`B�Ѕo � 0MGDI_�STA�%<q�! �� +0NC�c1\� ��
"~
"~d(/o�� �������#� 5�G�Y�k�}������� ŏ׏鏀% ��$�6� D�\qD�j�|������� ğ֟�����0�B� T�f�x���������ү L�����'�9�S�]� o���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ��������� �1�K�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�C�9� _�q������������� ��%7I[m ��������� !�M�Wi{� ������// //A/S/e/w/�/�/�/ �/���/??+?E O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�/�O �O_#_=?G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�O�o�o	5_ 'Qcu���� �����)�;�M� _�q����������oŏ ���-?I�[�m� �������ǟٟ��� �!�3�E�W�i�{��� ����ˏݏ����� 7�A�S�e�w������� ��ѿ�����+�=� O�a�sυϗϩ�#�կ ������/�9�K�]� o߁ߓߥ߷������� ���#�5�G�Y�k�}� ������������� '�1�C�U�g�y����� ����������	- ?Qcu����� ����;M _q������ �//%/7/I/[/m/ /�/�/���/�/�/ �/)3?E?W?i?{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O�/ �/�O�O�O_!?+_=_ O_a_s_�_�_�_�_�_ �_�_oo'o9oKo]o oo�o�o�o�O�o�o�o �o_#5GYk} �������� �1�C�U�g�y����� �o��ӏ����-� ?�Q�c�u��������� ϟ����)�;�M� _�q���������˯ݯ �	��%�7�I�[�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �������������� /�A�S�e�w߉ߛ߭� ����������+�=� O�a�s���ϱϻ��� ������'�9�K�]� o��������������� ��#5GYk} ������� 1CUgy�� �����	//-/ ?/Q/c/u/�/��/�/ �/�/��/?)?;?M? _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�/�/�O�O�O�O? _!_3_E_W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�O�O�o �o�o�o�O+= Oas����� ����'�9�K�]� o����o����ɏۏ�o ���#�5�G�Y�k�}� ������şן���� �1�C�U�g�y����� ����ӯ�߯	��-� ?�Q�c�u��������� Ͽ����)�;�M� _�qϋ�}ϧϹ���� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�ϕ� ������������� /�A�S�e�w������� ��������+= Oa������ ���'9K] o������� �/#/5/G/Y/k/� �/�/�/�/��/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcO}/kO�O�O�O �/�O�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[ouO� �$ENETM�ODE 1]�E��  
�@�@�a�D�o�`�|hRROR_PR_OG %�j%F��oy�eTABLE  �k�OCU�guw�bSEV_N�UM �b  ���a�p�a_A�UTO_ENB � �e�c�d_NON�q ^�k�a�r_  *��p��p%��p��p�p+�p�x�,��tFLTR��vHIS�s�A�`�{_ALM 1_�k� ��D�|@+-�ȏڏ����"�r1�_�r�p  �k��q�bg��`TCP_VER !�j�!�o2�$EXTL�OG_REQh�9�y��SIZ���STKߙ�u�~��TOL  �A{Dzp��A ��_BWDG��L�H���b1�DI6� `�EL��d�AM�STEP^�p��`���OP_DO��aF�ACTORY_T�UNh�dɩDR_?GRP 1a�iR��d 	b� ��`���������glrw��qŖ��J ���T��f�w�a� ���������Ϳ����<�'�`�Kυ@<���>gυ@
 Ifٓ�Ϲ�`�k���������	�C`}d�C��N<�B�y{D� �@UUT`��UT ߉�$� E׻� �߀��OH�cEP]��O���#M����KA��x�?�� ���:6:N��,�9-�4�x�
�) ��� m�-���!o�念b�e�3
{F�EATURE �b�EH��a�Handling�Tool ��B�English� Diction�ary��4D S�t��ard���A�nalog I/�O����gle S�hift��uto� Softwar�e Update��matic B�ackup��E�g�round Ed�it���Came�ra��F��Cnr�RndImJ��o�mmon cal�ib UI|��n�c��Monito�r��tr��Rel�iab��DHC�P����ata A�cquis����iagnosA����ocument �Viewe����u�al Check Safety��~��hanced��4��s` Frt���xt. DIO ���fiD�end.� Err��LC�J�s�	r���  7����FCTN Me�nuy v��*TPw Infac@��GigERd\��p Mask Ekxc� g�HTP�Proxy Sv�a�igh-Spe� Ski���< ~� mmunic@�7ons�ur7�	��Sconne�ct 2	(ncrRstru��*0 �eWq JC��KA�REL Cmd.� L�ua�g#R�un-Ti� Enyv](el +D��sB�S/W��Licenses`� �Book(Sys�tem)��MAC�ROs,�/Of'fse��%H� *��� MR����BMechStop�t  (�%i�	�\6ax� ��B�>od�witch�?037y.6�;Optm�?�03�fil`/7g���%ulti-T��f��PCM fun:'8Io%t1D^XMRegi� r�;FriY FHK�F��Num SelT5|�I�  Adju��N�A	��Mtatu��A�O[
��RDM �Robot��scgove��8Uea)@�� Freq An;ly�RemR0��n��8UDRServ�o� �0��SNPX� b�"�SNPC�liX�^
�Libr���_�� c4�P�V�o� t7ssag1E��{� �1��{��/IQ4eMILI�B]o7bP Fir�m(�GnP7Acc<]�e�TPTX5deln0zo8a�� 5�Hmorqu�imGula��z��fu�0�Pa�!Gn\���3&Χev.4e �ri�q �oUSB poort ��iP� �aY �vR EVN�Tw�pnexcept� yPfD�u���VC��r��X8V@$ ��o��[�S�PsSC�eH�SGE]��S�UI��Web PlV���Q������WZDT Appl���v����GridHQpla�y�D`I�&�R�r.���`�7�;R-20�00iC/125�L��2D Gui�pZ����Grap�hic����DV-� Path Ct�r��������dvn�DCS<pckw!���larm Caouse/wPed��Ascii��BL�oad` \�Upl�r��toS��%pr�ityAvoideM��l����Gu��P��¢8���s��t����yc��"�@rp~ ���5�os./�c�u �z��%	tr�ans.betw�.CRLmain �N��Q.��therNetZaz���`Ɵ�ca ��,RA�<p� ��(&0~Q/C�@o�'���L�<�o8�89���NRT����On��e Hel`��<E�@�AQ�tr�OROS ��7�e�⟨ ����sup�rt���vHap0A�[����Pk���GiG� t��Im��0F�0X�P�nsp� !+�|�64MB �DRAMdώ�FR�O�����l�ell����sh�����c��;��%�p>v�ty"�s�B��� r�B� �_R�0���~�3����hxP���MAIL⋞}�r �[�CP4�R��q�T1��[<��!Adp.G�X�As����/4Lz�CarHQq�Z�%Ro���+ax���OPT Pؿ�Ac'`��TX�!qpXpSyn.(�RSS)TVquir<`��DR�UT��^\� (�uess�S��h�]�V�RS6�duXp��[?��Pmi��3DLb�^�w!e��}K�`l Bui)@=n�APLCK�V�Հ�CGUxCRG���DD@��3LS���BU���1K�! /V�TAT*&�B��C*^�X/TCB@m/&4/~'x�~'F�/�&p~'�
7�u?TCEH1?C6�B7Vi?C6\�
6FP/�7l/
6�G�/�7�?�7?
6H,O
6IAIO[FHO
6LN�O+%MO�G�/H�G/
6N�O
6PdOHW�?
6R�?
6SD_rW`_
6W�_�W_
4gVGF�_�UP2� �W�O�W�_�VB@o�V	D\o�VF�/�VO�7TUT<b01�o�fy2�o�bTBGG$br�lr~��� UI�`�|�HMI"r�po�n��`�Q�for �s�>s�KARELK��al�TPY�c|��|������� ���*�<�i�`�r� ������Տ̏ޏ�� �&�8�e�\�n����� ��џȟڟ����"� 4�a�X�j�������ͯ į֯�����0�]� T�f�������ɿ��ҿ ������,�Y�P�b� �φϘ��ϼ������� ��(�U�L�^ߋ߂� ���߸������� �� $�Q�H�Z��~��� ����������� �M� D�V���z��������� ������
I@R v������ �E<N{r �������/ /A/8/J/w/n/�/�/ �/�/�/�/�/�/?=? 4?F?s?j?|?�?�?�? �?�?�?�?O9O0OBO oOfOxO�O�O�O�O�O �O�O_5_,_>_k_b_ t_�_�_�_�_�_�_�_ o1o(o:ogo^opo�o �o�o�o�o�o�o - $6cZl��� �����)� �2� _�V�h�������ˏ ԏ���%��.�[�R� d�������ǟ��П� ��!��*�W�N�`��� ����ï��̯ޯ�� �&�S�J�\������� ����ȿڿ���"� O�F�Xυ�|ώϻϲ� ���������K�B� T߁�xߊ߷߮����� �����G�>�P�}� t���������� ��C�:�L�y�p��� ����������	  ?6Hul~�� ����;2 Dqhz���� �/�
/7/./@/m/ d/v/�/�/�/�/�/�/ �/?3?*?<?i?`?r? �?�?�?�?�?�?�?O /O&O8OeO\OnO�O�O �O�O�O�O�O�O+_"_ 4_a_X_j_�_�_�_�_ �_�_�_�_'oo0o]o�Tol  �H552oc�a21n�eR78�h50�e�J614�eATU]P�f545�h6�e�VCAM�eCRIn�gUIF�g28�f�NRE�f52�fR�63�gSCH�eDwOCVOvCSU�f�869�g0�fEI�OC+w4�fR69��fESET�g�gJ�7�gR68�fMA{SK�ePRXYx]7�fOCO�x3�hh�f�p�h3�vJ6�h�53rvH$�LCH^�vOPLG�g0��MHCR�vSm�MkCS�h0�w55�f�MDSW���OP��MPR�?p2�0n�fPCMvR0����p�fw�2�51�g5u1.�0�fPRS�w�69�vFRD�fFwREQ�fMCN�f{93�fSNBA7w^%�SHLB��M��t?p��2�fHTC�f�TMIL�hrvTP�A�vTPTX�EL��w�rw8�g�`�fwJ95vTUT��95�vUEV�vU�EC�vUFR�fV�CC��O��VIP���CSC�CSGt*vdpI�eWEB�f7HTT�fR65x@��CG��IGݧIP�GS�RC��DG��H72�w9Q�R76�fR8��w�b�;85rvR66b��w�R,�R51�w53�"�68n�66�2��6.�6vJ74�g75b���`b�<��R5Y�J59.�5�8.�85�54��6nm�NVD�vR6y�,���87j�4v�p�:�i�R7w�pvDu0m�F�RTS���CLI��gCMS��v?��fSTY��6���CTO�fcp�w7�qxNN
�NN�vO�RS���pF�3��5�HPM�z�\�?p��fOPI2�3�ڸ7�rvCPR��L��S���7�vSVSNvS;LM�vV3D��wwPBV�APL�vwAPV�CCG�f�CCRn�CD��C�DL2�CSBfvC�SKCT�CT1Bަ�TC�����CҧTCv���TC��TC�vCT1ENvs��TEZvs�VƧTF
�F�G��G��^�H^�I�Tv�CT)�CTM���� ��N^�P��P���R
�A�TS
�W�r	2�VGF�P2F��P2��� �B��D�FvV�VT��g� �fVTB��V�ewIH�V;�K��V��vhQcu� ������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?m??�?�?�?�? �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_e_w_ �_�_�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9K]o���� �����#�5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�W� i�{ߍߟ߱������� ����/�A�S�e�w��  H5�5y�����R7�8��50��J61�4��ATU����5�45��6��VCAܢ��CRI�UI����28�NREv��52�R63���SCH��DOCVr��C��869��0��EIO2e�4��R69�ESE�T���J7�R6�8��MASK��P�RXY?�7��OC�O3��� ��3�n
J6��53��H�LCHN
OPL�G��0�
MHCR�O
SMCS��0�55��MDSW�o}OP}MPR�~
{�0��PCM>�R0� ���[51��51,0��PRS69n
F{RD.�FREQ��MCN��93��S�NBAo��SHLEB�*M�+{�^2���HTC��TMILܯ��TPA��TPTX:EL�*��q8���~�J95N��TUT~95n
U�EV
UECN
U�FR.�VCC�<O�.VIP:CSCNN:CSG^���I��wWEB��HTT��R6m�|<CGmKI�GMKIPGS�JR�C:DG}H72���9=+R76��R�8]P�K85��R�66�L��R,R5m1��53�68[�66�2�6,6nN�J74��75�L�����K�R5�;J[59k58k8m<�54n[6[NVD�
R6[P�87�^l4N�; l]+R7XM�; N�D0[F,|wRTS�*CLI����CMS��{p��S�TY;6mCTOh�����7��NN�[;NNn
ORS.; �.l3�k5�[HPM�L,{���OPI�Jkp�\7��CPR�~+L�;S�7n
S�VS��SLM
Vs3DL=�PBVN:wAPL��APV~
wCCG��CCR�CD�;CDL�JC�SB��CSK~CT=;CTBNJېK�TC�*��ΜC>KT�C>���^�TC��TC
CTE��k�n�cTE��k�.KTFޜ�F�GΜG��N�HjN�IN{T��CT];�CTM�M�;���N*N�P�PΜRޜ}|�TSޜW���JVGmF޻P2�;P2�*T���B�D�F>��V��VT��k���VkTB~�V��IH;)V�@��KKVmJ~� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi{���� ���/AS ew������ �//+/=/O/a/s/ �/�/�/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� �������� %�7�I�[�m������ ��Ǐُ����!�3� E�W�i�{�������ß ՟�����/�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�� �'�9�K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}ߏߡ߳� ����������1�C��U�g�y���S�TD��LANG������������ �"�4�F�X�j�|��� ������������ 0BTfx��� ����,> Pbt����� ��//(/:/L/^/ p/�/�/�/�/�/�/�/� ??$?6?H4RBT��OPTN_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O�O�O�O�ODPN��	__-_?_Q_c_ u_�_�_�_�_�_�_�_ oo)o;oMo_oqo�o �o�o�o�o�o�o %7I[m�� ������!�3� E�W�i�{�������Ï Տ�����/�A�z� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7opIo[omod99{e��$FEAT_A�DD ?	�����a�`  	zh�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������# 5GYk}��� ����//1/C/�U/g/y/�/�/�dDE�MO b�i   zh�-�/�/ ??"?O?F?X?�?|? �?�?�?�?�?�?OO OKOBOTO�OxO�O�O �O�O�O�O___G_ >_P_}_t_�_�_�_�_ �_�_oooCo:oLo yopo�o�o�o�o�o�o 	 ?6Hul ~������� �;�2�D�q�h�z��� ��ˏԏ���
�7� .�@�m�d�v�����ǟ ��П�����3�*�<� i�`�r�����ï��̯ ����/�&�8�e�\� n���������ȿ��� ��+�"�4�a�X�jτ� �ϻϲ���������'� �0�]�T�f߀ߊ߷� ����������#��,� Y�P�b�|����� ��������(�U�L� ^�x������������� ��$QHZt ~������  MDVpz� �����/
// I/@/R/l/v/�/�/�/ �/�/�/???E?<? N?h?r?�?�?�?�?�? �?OOOAO8OJOdO nO�O�O�O�O�O�O_ �O_=_4_F_`_j_�_ �_�_�_�_�_o�_o 9o0oBo\ofo�o�o�o �o�o�o�o�o5, >Xb����� ����1�(�:�T� ^�����������ʏ�� � �-�$�6�P�Z��� ~�������Ɵ���� )� �2�L�V���z��� ����¯����%�� .�H�R��v������� ������!��*�D� N�{�rτϱϨϺ��� ������&�@�J�w� n߀߭ߤ߶������� ��"�<�F�s�j�|� ������������ �8�B�o�f�x����� ��������4 >kbt���� ��0:g ^p������ 	/ //,/6/c/Z/l/ �/�/�/�/�/�/?�/ ?(?2?_?V?h?�?�? �?�?�?�?O�?
O$O .O[OROdO�O�O�O�O �O�O�O�O_ _*_W_ N_`_�_�_�_�_�_�_ �_�_oo&oSoJo\o �o�o�o�o�o�o�o�o �o"OFX�| �������� �K�B�T���x����� ����������G� >�P�}�t��������� ������C�:�L� y�p����������ܯ ���?�6�H�u�l� ~��������ؿ�� �;�2�D�q�h�zϧ� �ϰ������� �
�7� .�@�m�d�vߣߚ߬� ���������3�*�<� i�`�r�������� �����/�&�8�e�\� n��������������� ��+"4aXj� �������' 0]Tf��� �����#//,/ Y/P/b/�/�/�/�/�/ �/�/�/??(?U?L? ^?�?�?�?�?�?�?�? �?OO$OQOHOZO�O ~O�O�O�O�O�O�O_ _ _M_D_V_�_z_�_ �_�_�_�_�_o
oo Io@oRoovo�o�o�o �o�o�oE< N{r����� ����A�8�J�w� n���������Џڏ� ���=�4�F�s�j�|� ������̟֟���� 9�0�B�o�f�x�����>ȭ  ��ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ �������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/�/�/�/�)  �(�!�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |������� ��0�B�T�f�x��� ������ҏ����� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� \�n������������� ����"4FXj |������� 0BTfx� ������// ,/>/P/b/t/�/�/�/�/�!� �(�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFoXo jo|o�o�o�o�o�o�o �o0BTfx �������� �,�>�P�b�t����� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�D�V�h� z�������¿Կ��� 
��.�@�R�d�vψ� �ϬϾ��������� *�<�N�`�r߄ߖߨ� ����������&�8� J�\�n������� �������"�4�F�X� j�|������������� ��0BTfx ������� ,>Pbt�� �����//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? �?�?O O2ODOVOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����������Ω�$FEA�T_DEMOIN�  Ӥ�����Ԡ�INDEX�����ILE�COMP cw���4����*�SETUP2� d4�>���  N i�'�_�AP2BCK 1�e4�  �)�Ϩ����%��пԠ 7�����ѥ��'϶�K� ڿXρ�ϥ�4����� j��ώ�#�5���Y��� }ߏ�߳�B���f��� ��1���U�g��ߋ� ����P���t�	�� ��?���c���p���(� ��L���������; M��q ��6� Z�~�%�I� m�2��h ��!/3/�W/�{/ 
/�/�/@/�/d/�/? �//?�/S?e?�/�?? �?�?N?�?r?O�?O =O�?aO�?�O�O&O�O JO�O�O�O_�O9_K_ �Oo_�O�_"_�_�_C��w�P{� 2���*.VR�_o�P*oCo�SIomoWU`�PCuo�o�PFR6:�o�nYo�o}kT�$�eN|��x�otVV*.FoD��Q	�c��|a��{STM�+��b��`�V��z��{H G���<���X�j����zGIF	�3�>��܏8��zJPG�����>���`�r��~jJS��:��P͓(��%�
JavaScrgiptf���CSW��=���h� %C�ascading� Style S�heets�\P
�ARGNAME.SDT�|\A�\-���M�]�n��]�DISP*d�G�A����񿀵�򿞿
TP�EINS.XML�!�Ϳ:\5��U�C�ustom To�olbarvϥ�PASSWORD�~z^FRS:\���x� %Pass�word Con�fig�Ϧ���� Y�@���ϥ�W_��{_ ���߱_#��G�Y��� }����B���f��� ����1���U���y��� ���>�����t�	�� -?��c���� �L�p�; �_q �$�� Z�~/�/I/� m/��/�/2/�/V/�/ �/�/!?�/E?W?�/{? 
?�?.?�?�?d?�?�? O/O�?SO�?wO�OO �O<O�O�OrO_�O+_ �O$_a_�O�__�_�_ J_�_n_oo�_9o�_ ]ooo�_�o"o�oFo�o �o|o�o5G�ok �o��0�T�� ���C��<�y�� ��,���ӏb������ -���Q���u������ :�ϟ^�ȟ���)��� M�_�������H� ݯl�����7�Ư[� �T��� ���D�ٿ� z�Ϟ�3�E�Կi��� �ϟ�.���R���v��� ߬�A���e�w�ߛ� *߿���`��߄��+� ��O���s��l��8� ��\������'���K��]��������� ��$FILE_DG�BCK 1e�������� < �)
S�UMMARY.DyG��e�MD:���-q�Diag� Summary�.;�
CONSLOG#q�@�Console� log�:�	T�PACCN�%��1<TP A�ccountin��;�FR6:I�PKDMP.ZI	Pei�
}�=M�Exceptio�n�;�*.DT��/q�FR:\��>.�FR DT Files>/�j MEMCHECCK'��/��Memory D�ata�/��(i{\)�!RIPE�p�/�/A?�#%1� Packet 9L��%�b"1STAT;?"?4?�?� %]2St�atu_/y<	FTAP?!O�?%O�'��mment TB�DNO�'��)ETHERNE�?�&O�!�O�O@Et�hernf0� fi�gura�A�8ADCSVRFBO(O:O�S_�3P verify allV_��$���UDIF�FK_1_C_�_W3mXd�iff�_�W�!PCHG01�_�_�_]o��1�_�o�R�i2 So:oLo�o�_�o�o"b�3�o�o�oe ��o�vVTRNDIAG.LS��BT��!�q O�pe�Ch1 Eno�stic�'�<�)VDEV�rD�A0/��m��1V�is�Devic9e� �IMG�r��H�Z��V3��Imsag���UP6��ES5�ʏFRS�:\5�@/B Upd�ates Lis�tv�;�݀FLEXEVEN�OΏ������1�� UIF� EviAi?�#����)
PSRBW�LD.CM%�e��a�=�x�� PS_R?OBOWELoO9��AIOׯ����'��BNet/IP�pa"��#ߌ)��GRAPHICS4D������%4D Gr?aphicsZ/�'w�' 2GIG?��o���&GigqE���#���2�SMOc����'~P�/Email$��=��\��SHAD�OW��h�z���#�Shadow C�hang���& �~��RCMERR�����ϓ��#X�CFG Error���t��6� �+���3CMSGLIB ��r߄������2��x�����*�)��ZDT�s����'�ZD0�ad9���&=쿢NOTI_v������%Noti�fic�B���&�A�)��u�X�d������������������� ��AS��w� *<�`��+ �O�H��8 ��n/�'/�� ]/��/�/"/�/F/�/ j/�/?�/5?�/Y?k? �/�??�?B?T?�?x? OO�?CO�?gO�?`O �O,O�OPO�O�O�O_ �O?_�O�Ou__�_�_ :_�_^_�_�_�_)o�_ Mo�_qo�oo�o6o�o Zolo�o%7�o[ �ox�D�h ���3��W��� �����ÏR��v�� ���A�Џe�􏉟�� *���N��r������ =�O�ޟs����&��� ͯ\�񯀯�'���K� گo������4�ɿۿ j�����#ϲ��Y�� }�ϡϳ�B���f��� �Ϝ�1���U�g��ϋ� ߯�>ߨ���t�	�� -�?���c��߇��(����x��$FILE�_FRSPRT � ����������MDONLY 1e���|� 
 �)�MD:_VDA�EXTP.ZZZ���z�Q�`�6%�NO Back? file +�B��U�W��A��� ����Q�0��Tf �����O�s �>�b�o �'�K���/ �:/L/�p/��/�/ 5/�/Y/�/}/�/$?�/ H?�/l?~??�?1?�?��?g?�?�? O2O��VISBCK	����*.VD3O}O�0�FR:\L@ION\DATA\hO��2�0Vision VD~�O�8?*.CAM�O_� %	�A�C�O�L�GigE Cam�era Definit�@-_�?}_�? �_O�_�_f_�_�_o 1o�_Uo�_yo�oo�o >o�o�oto	�o-�o &c�o���L �p���;��_� q� ���$���H���� ~����$�I�؏m�7N�LUI_CONF�IG f��|_A|� $ Z��{��ӟ���	��-�;���|xc�e�w� ��������S���� �(���9�^�p����� ��=�ʿܿ� ��$� ��H�Z�l�~ϐϢ�9� ��������� ߷�D� V�h�zߌߞ�5����� ����
���@�R�d� v���1�������� ����<�N�`�r��� ������������� &8J\n�� ������"4 FXj|��� ����/0/B/T/ f/x//�/�/�/�/�/ �/�/?,?>?P?b?t? ?�?�?�?�?�?w?�? O(O:OLO^O�?�O�O �O�O�O�OsO __$_ 6_H_Z_�O~_�_�_�_ �_�_o_�_o o2oDo Vo�_zo�o�o�o�o�o ko�o
.@R�o v�����g� ��*�<��M�r��� ������Q�ޏ���� &�8�Ϗ\�n������� ��M�ڟ����"�4� ˟X�j�|�������I� ֯�����0�ǯT��f�x�������A�R�obot Spe?ed 10%��鿠����1�?�H�x�8�E��$FLUI�_DATA g����u��?�g�RESU_LT 2hu���� �T�/�wizard/g�uided/st�eps/ExpertT��������߀/�A�S�e�w߉ߗ��Skip G���ance and� Finish Setup������ ���"�4�F�X�j�|�\��<� H�.?��uŷ�0 ��H�����u����ps��"�4�F�X�j�|� ��������������H� !3EWi{� �����?���?������+��&��ri�p����ToolN�um/NewFrame����� ���//*/</��0x0?/g/y/�/ �/�/�/�/�/�/	??-???  <�;�?����dime?US/DSTB?�? �?�?OO/OAOSOeO�wO�O��Enablv�O�O�O�O__�)_;_M___q_�_�_F�G��?q?�_�?�?�224�?%o7oIo[o moo�o�o�o�o�o�O �O!3EWi{ �������_�_p�_,��_ ozon�0 �}�������ŏ׏������1���ES�T Ea��rn St�Э�;�t����� ����Ο�����(�X:���J� �?�7���{���Ϻ�Region>�ͯ߯�� �'�9�K�]�o������America ���Ϳ߿���'π9�K�]�oρ�@�R�y��i����ϟ�bEditor��!�3�E� W�i�{ߍߟ߱����������ular �
�� (reco/mmen�)��(� :�L�^�p���������G�������#������/acces ��t����������������(?�Co�nnect to� Network 7n������@��"4K�����s��!I�_�I�ntroduct �����//&/8/ J/\/n/�/C�p�/�/ �/�/�/�/??0?B? T?f?x?�?�rR��r��i�?9��/Safet��O O2ODOVO hOzO�O�O�O�O�O�/ �O
__._@_R_d_v_ �_�_�_�_�_�_�?�? �_'o�?W�j�oo�o�o �o�o�o�o�o�o# �OGYk}��� ������1��_�oov�8i#EoWf/current8� ͏ߏ���'�9�K��]�o���D15-M�AY-20 09?:31 AM���� П�����*�<�N�`�r������烏e��ǯ5l ����Yea ��/�A�S�e�w����������ѿ@2020ۿ��(�:�L� ^�pςϔϦϸ������ 
����  �෯ߋ��Month��s߅ߗߩ߻߀��������'�B5/�U�g�y���� ��������	��-���F�� �m�3nA���DaO�������� 0BTfx��1C����� '9K]o�@�R�_��ۯ����Hou�/+/=/O/ a/s/�/�/�/�/�/8�9�/�/?!?3?E?W? i?{?�?�?�?�?�?�"R�	�O3n"�S�inute�?pO�O �O�O�O�O�O�O __$_�31+_R_d_v_ �_�_�_�_�_�_�_oo*o�?S�Oio�=O��AMP���o�o �o�o	-?Qc u�������� ��"�4�F�X�j�|�*����攠{o]o俏-L�o��NetDon^O�#�5�G� Y�k�}�������ş� Z������1�C�U� g�y���������ӯ8aACo����;�&冿ripperO�o�olNum/FraX�s �o������� ��ɿۿ����#�>� @_L�^�pςϔϦϸ� ������ ��$�;oQ�����i�/J)9�K�ActiveW�*��� �������!�3�E�W�<i�(�0x0{�� �����������!�3�pE�W�i�{�  =���������ߗ�MacSroS���w��s~� -?Qcu�� ��|���) ;M_q����@�������/.K,��<����Open\�o/ �/�/�/�/�/�/�/�/ ?�:�G?Y?k?}?�? �?�?�?�?�?�?OO�6�H�/dO֏�Summary&O�O�O �O�O�O_"_4_F_X_ j_ٟ�_�_�_�_�_�_ �_oo0oBoTofoxo���[O�oO�RobotOp|o
 .@Rdv��� �}_����*�<� N�`�r���������̏ �o�o�o��f-5/G/oClos[�k�}� ������şן�����2�E�W�i�{� ������ïկ������4OFI��]��n�1��BetMethod"���ǿٿ�����!�3�E�W�i�,7�Direct e�ntry of �EOAT datasϱ����������@�/�A�S�e�v��@]�RB�U����h$����Btraight?Offsetv��  �2�D�V�h�z�������12�� Tool������/�A� S�e�w���������~� ��ߤ��m%�ߚA��AX��cu�� �����21�298.499 3�GYk}���@����/-5�C�?���]/1CY/�/�/�/�/ �/?#?5?G?Y?k?�q�	-169.1565o?�?�?�?�?�? �?	OO-O?OQOcO"/<4/���)(O/�Os/�/CZrO__/_ A_S_e_w_�_�_�_�_�*951.8884�_�_oo&o8oJo \ono�o�o�o�ouO�O�CDm�ۣO���)�O��Rotation=wW�ocu ����������_179.868�?C�U�g�y����� ����ӏ���	��o�oD%3�V�oY�-?P���ɟ۟�����#�5�G�Y��-.2586k����� ��̯ޯ���&�8��J�\��-�g���hAK���o�����Rn� ��/�A�S�e�wω���ϭ�l�-29.4700������� "�4�F�X�j�|ߎߠ���q�������ȟ���J"ѿ�tp�3Zdir/Tp3z��X�j�|��� ������������_0� B�T�f�x��������� �����������o��_Ͱ+%��Mea�surement�/Straigh �O����� 1CU�&���� ����	//-/?/ Q/c/"4F�/j|�/We�Nums//New�#sj/	? ?-???Q?c?u?�?�?�?j0x���?�? OO*O<ONO`OrO�O�O�O�Op}/�I�/��O�.�/�,Tool�#Use�O`_r_ �_�_�_�_�_�_�_om1o5oGoYoko }o�o�o�o�o�o�o�oDp
�OQp�O�M_!_�,Part F_������� )�;�M�_�b2c��� ������я�����@+�=�O�a� 2y?䡟�(u�'s/G ڰ�#f���&�8�J��\�n����������71.10���� ��)�;�M�_�q����������|/�&B�3�3�����)ɟۙP�ayload1Cm�V�h�zόϞϰ����������
��E�OAT with tot�=�O�a� s߅ߗߩ߻��������oͿ�O)�S��� 'ϔy������������(�:�L�^��.Ϡѯ���������� ����*<N`˿1z ?��u�3�2C�� 2DV@hz���Ǡ�no(���//'/ 9/K/]/o/�/�/�/� v4��/�/ns&��	�Advanced �/P?b?t?�?�?�?�?��?�?�?OǠ0x w�.O@OROdOvO�O�O��O�O�O�O�O_�� �/�/%_O_mt%?��Mass/Center�Q
_�_�_�_ �_�_�_o!o3oEoWo~ơ-32.3u� �o�o�o�o�o�o�o�'9K]tڶ�鿛�o_�^��^ ���1�C�U�g�y�����\onb2toُ� ���!�3�E�W�i�{��������p�w ��H��z,��G"0	c�R�xX��R�d�v� ��������Я���c�1.5ȏ+�=�O� a�s���������Ϳ߿0�� �?��C���)��RYϦϸ� ������ ��$�6�H�~�-.1999W� �ߔߦ߸������� ��$�6�H���Sž�Lៗ�Y�k�}ύRZ Z�����0�B�T�f� x�������qo������ ,>Pbt����i�����x.����p�p�|@�Oa s������� ���'/9/K/]/o/�/ �/�/�/�/�/�/�/��(��D?*rt �ϣ?�?�?�?�?�?O !O3OEO\�n�{O�O�O �O�O�O�O�O__/_ A_S_?|�6?�_Z?l?~?rt���_	oo-o ?oQocouo�o�o��Ə �o�o�o);M _q���f_ԟ�_�����\TCPVe�rify/&�Method�J�\�n� ��������ȏڏ쏫l�Direct Entry��,�>� P�b�t���������Ο���x���=�2�z'��fy>�� ����ί����(��:�L���298.4992O�|������� Ŀֿ�����0�B�x��M�C�?�/� ��S�e�#��?����� "�4�F�X�j�|ߎߠ����	-169.1565��������� �+�=�O�a�s���xV�h�&2�)(�� ��Ϲ�#��_@�R�d� v�����������������a951.8884��$6HZl~ �����������Dm����9���#�W����� ��//%/7/I/�`179.868�� w/�/�/�/�/�/�/�/�??+?=?�x�3��V+�?Oa#�P N?�?�?OO1OCOUO�gOyO�O�O �-.2586�O�O�O �O __$_6_H_Z_l_�~_�_O?a?�5��hA?�_�?�?#�R�_ =oOoaoso�o�o�o�o��o�o�o`�-29.4700�o 2D Vhz��������_�_�S����_5��Z*oofyMean������� ʏ܏� ��$�6��o*[�G�t��������� Ο�����(�:�� �i�'����Z)Y�k�}�axJ������ /�A�S�e�w���H�Z� ��ѿ�����+�=� O�a�sυϗ�V���z�����["����Int�roductio ��3�E�W�i�{ߍߟ� �������ߪE���� (�:�L�^�p���� ���������������9��R�tut�ojog��Overview����� ����������& 8��\n���� ����"4F���a���]�Se�lectT1ModeH�� //$/ 6/H/Z/l/~/�/O�/ �/�/�/�/? ?2?D? V?h?z?�?K]o�?��?`(���Ena�bleTeachPendant�? 6OHOZOlO~O�O�O�O �O�O�O�/_ _2_D_ V_h_z_�_�_�_�_�_@�_�?�?�?+oI�$�?^�Joinl`g�_ �o�o�o�o�o�o�o (:�O^p�� ����� ��$��6��_oo{����'|Qog�ride_mo Տ�����/�A�S� e�w���H����џ� ����+�=�O�a�s� ����V�h���ܯ��`��HoldDead�manSwitch��1�C�U�g�y��� ������ӿ忤�	�� -�?�Q�c�uχϙϫ� �����Ϡ�ίį&��=� ���ResetAlarm��~ߐ� �ߴ���������� � 2��V�h�z���� ��������
��.�@�A���[����!M��ą_J1@����� ��	-?Qcu �F����� );M_q����T�f���Lo��J2-J6�*/</N/`/ r/�/�/�/�/�/�/� ??&?8?J?\?n?�? �?�?�?�?�?����O1O�#�cgCarȏyO�O�O�O�O�O �O�O	__-_�/Q_c_ u_�_�_�_�_�_�_�_ oo)o;o�?OVo�o�&IO��eO�o�o�o '9K]o� @_������� #�5�G�Y�k�}���No`o��ԏ��o[A�d_X��!�3�E�W�i� {�������ß՟��� ��/�A�S�e�w��� ������ѯ㯢�����x(�����_Y-Z� w���������ѿ��� ��+��O�a�sυ� �ϩϻ��������� '����
�T�~�����_Rotation���������'� 9�K�]�o��@ϥ�� ���������#�5�G� Y�k�}�<�N�`߂����o��onc�!3E Wi{����� ���/ASe w���������8����(/�� ��[A�LastScreen�r/�/�/�/�/ �/�/�/??&?�J? \?n?�?�?�?�?�?�? �?�?O"O��/OO�yO;+file/b�ackup�ddevice4O�O�O�O �O_ _2_D_V_h_z_�96Front �Panel USB (UD1)�_ �_�_�_�_oo)o;opMo_oqo�o  EBA�CAOaO�o��%�O��Firectories�o1CU gy�����>1��P:\\BKU�P_12-DEC�-18_01-4?8-30\\�� -�?�Q�c�u������� ��Ϗ�mJO�o�o$�B��oE�defڏo��� ������ɟ۟�����#�:5Image B�B+�\�n����� ����ȯگ����"��m�=@'�	�k����A%gripp�erP$ToolNum.���ѿ���� �+�=�O�a�s�6?�� �ϻ���������'� 9�K�]�o߁�DOR�d��������S!G��Typ�O�%�7�I�[�m��������Single �� ������*�<�N�`��r������������lg��o��!�g��Co�mment/cmt��o�����@���#���� L^p�����@�� //$/�����#g/-�?���Summary*/�/�/ �/�/??+?=?O?a? s?�ϗ?�?�?�?�?�? OO'O9OKO]OoO�� @/R/�O�O�!"�/�eprogres _%_7_I_[_m__�_ �_�_�_�?�_�_o!o 3oEoWoio{o�o�o�o�o�m�O�O�o�",�O�M�F6�or� ���������\-#�I�[�m�� ������Ǐُ���� !�8/�of�(:Lss7&�Ɵ؟����� �2�D�V�h�'�0 w�������ӯ���	� �-�?�Q�c�u�4�F��X���|�����ss8 z��,�>�P�b�tφ��Ϫϼ��\Ini�tializ�� B�"����'�9�K� ]�o߁ߓߥ߷��߈�������,	9KIO/s1��a�s�� ������������ ,�O�D�V�h�z����� ����������
�B
���A��]�1�C�2"����� !3EWi(�� ������//�(/:/L/^/p//A
�O�/�N!��Commentv/?? /?A?S?e?w?�?�?�? �?�_�?�?OO+O=O OOaOsO�O�O�O�O�MA�/���O_�/ � �OS_e_w_�_�_�_ �_�_�_�_oo�?=o Ooaoso�o�o�o�o�o �o�o#g�O�O ;e.o���� ����!�3�E�W� i�(o������ÏՏ� ����/�A�S�e�v�JpkE����{�� ���(�:�L�^�p� ��������w�ܯ� � �$�6�H�Z�l�~��� ����s��������͟ 2�D�V�h�zόϞϰ� ��������
�ɯ.�@� R�d�v߈ߚ߬߾��� ������׿���]� τ���������� ��&�8�J�\�߀� �������������� "4FXj)�;�M���(-_�!MacroNumA_  $6HZl~�� �s����/ /2/ D/V/h/z/�/�/�/�/ �O��/?�!���easurement�/W?i?{?�?�? �?�?�?�?�?O�/O AOSOeOwO�O�O�O�O �O�O�O_�/�/�/4_�^_� %?71Weight��_�_�_�_ �_ oo$o6oHoZoO ~o�o�o�o�o�o�o�o  2DVh'_9_K_��y_�W�_� ��0�B�T�f�x��� ����moҏ����� ,�>�P�b�t������� ��{���s�(�:� L�^�p���������ʯ ܯ� ���$�6�H�Z� l�~�������ƿؿ� ���}ߟ�S��z� �Ϟϰ���������
� �.�@�R��c߈ߚ� �߾���������*� <�N�`�ρ�Cϥ�g� ��������&�8�J� \�n������������� ����"4FXj |���q����� ��0BTfx� ������/�� ,/>/P/b/t/�/�/�/ �/�/�/�/?�%?� I??�?�?�?�?�? �?�? OO$O6OHOZO /~O�O�O�O�O�O�O �O_ _2_D_V_?w_ 9?�_�_qO�_�_�_
o o.o@oRodovo�o�o �okO�o�o�o* <N`r���g_ �_�_���_&�8�J� \�n���������ȏڏ ����o"�4�F�X�j� |�������ğ֟��� ���'�Q��x��� ������ү����� ,�>�P��t������� ��ο����(�:� L���/�A���e��� ���� ��$�6�H�Z� l�~ߐߢ�a������� ��� �2�D�V�h�z� ����oρϓ���� �.�@�R�d�v����� ������������* <N`r���� ���������G 	�n������ ��/"/4/F/W/ |/�/�/�/�/�/�/�/ ??0?B?T?u?7 �?[�?�?�?�?OO ,O>OPObOtO�O�O�O �?�O�O�O__(_:_ L_^_p_�_�_�_e?�_ �?�_�?o$o6oHoZo lo~o�o�o�o�o�o�o �o�O 2DVhz ��������_ ��_=��_�v����� ����Џ����*� <�N�r��������� ̟ޟ���&�8�J��	�k�-������/�wizard/g�ripper/s�teps/SummaryU����� �/�A�S�e�w����� Z���ѿ�����+π=�O�a�sυϗϩ� � _�������W����ˡTCPVerifկ<�N�`�r߄� �ߨߺ������߯�� &�8�J�\�n���� ���������������C�]�"�ˡG IO&ߎ����������� ��0B�fx ������� ,>PW �%� o�_�����/ /,/>/P/b/t/�/�/ W�/�/�/�/??(? :?L?^?p?�?�?W�i�w��?�O"O4O FOXOjO|O�O�O�O�O �O�O�/__0_B_T_ f_x_�_�_�_�_�_�_ �_�?�?�?;o�?boto �o�o�o�o�o�o�o (:�OKp�� ����� ��$� 6�H�oi�+o��Oo�� Ə؏���� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v�����Y���}�߯�� ��*�<�N�`�r��� ������̿޿𿯟� &�8�J�\�nπϒϤ� �������ϫ��ϯ1� ���j�|ߎߠ߲��� ��������0�B�� f�x���������� ����,�>���_�!� ����Y�������� (:L^p�� S���� $ 6HZl~�O��� s�����/ /2/D/ V/h/z/�/�/�/�/�/ �/�
??.?@?R?d? v?�?�?�?�?�?�?� ��O9O�`OrO�O �O�O�O�O�O�O__ &_8_�/\_n_�_�_�_ �_�_�_�_�_o"o4o��?OO)O�oIC�$�FMR2_GRP� 1i�e�� �C4 w B�KP	 KP��o�l�`E�� ��o�G[�`OHcE�P]��O��#�M��-qKA���}?pIEl�`:6:N�uq�9-�}u}A��  ��{BH�cC`}dC��N�qOB�{�uEl�dx���`@UUT��UT}�R��a>F�D�>�d�>D��=�=��1U�op�H$:���=:��:�.�	:sf�:�Uf1���}������ۏ���8�KW�b_C�FG j�kT �C�������J�N�O �jF�236039 9�737K�RM_C�HKTYP  ��aKP�`�`�`�aRO=M��_MIN��KSW��+���pX�`�SSBZ�k�e �fX�KU�O�x���P�TP_D�EF_OW  �KT�c��IRCO�M�����$GENOVRD_DO ��VQݭTHR � �d��d�_ENB�ϯ �RAVC�clA�L� ���f��`�}E����G
�F�?/lG�,�t�4��KR�`!��bv���r��C�kOU�`r�l KPq�h���e<(��[5�ۿ-�^������������]�^��<�,!�������n"���C����'c>D�j�pKQC�����W������B�`��B���a���i ɑ�D�SMT�csQ��`N�����$HAPTIC_CNT 2t�e�[�
!���@�W�KSs<x�A��KS��x�Cv�s2x�I�KS}���H���s�^@x�E�Ԗ����ȹKS�6x�Gɺ��KPZ�pz�q�͐KS!�Z�FE�AT  g�Z�� <�8��B�T�c��X�OST_�\�1uܴiM��V_ 	�������KV��HYe���$�6� H�HZ �y������������f�	anonymous��(:L ������ ��h���Z�7 I[m������ ���/Vhz� �{/��/�/�/�/�/ .??/?A?S?v/� ��?�?�?�?�?*/</ N/+Ob?OO�/sO�O�O �O�/�O�O�O__8O 9_�?]_o_�_�_�_�? �?O"O$_�_XO5oGo Yoko}o�O�o�o�o�o �ooB_T_1CUg y�_�_�_��o�,o 	��-�?�Q��u��� �����Ϗ��� )�;�������̏ �˟ݟ���Z�7� I�[�m����؏�ǯ ٯ����V�h�z��� ��{�����ÿտ� .���/�A�d�RϬ���ϛϭϿ����w�E�b�1v���  CP!e�#����� N�=�r�5ߖ�Yߺ�}� �ߡ������8���\� ��C��g�y���� ����"���F�	��|� ?���c����������� Bf)�M �q����, �Pt7I�m�����QUI�CC0��!1?1.200.@!&/r)1O/+/!  @/�R/!2�/{/��/!ROUTER�/��/!
?$� ?��PCJOG???�!192.16�8510�/#CAMgPRT�?k?!511�0�?�6RT?�?��?-O��NAME �! �!ROB�O�?5OS_CFG� 1u � ��Auto-started6�/FTPA��AX� Z��O��_'_9_K_]_ ���_�_�_�_�O�_n_ �_o#o5oGo��O�O �O�o�_�O�o�o�o �_BTfx��o /������� 1�C�U�����o���� Ώ����(�:�L� ^����������ʟܟ �5�G�Y�6�m�Z��� ~�������{�د��� � �C�ů?�h�z��� ������	��-�/�� c�@�R�d�vψ�O��� ��������ϙ�*�<� N�`�r߄�˿ݿ��� ���7��&�8�J�� ���������m� ���"�4�F��ߟ߱� ������������� ��BTfx��� /����a� s���3������ ����/(/:/L/ op//�/�/�/�/�/�pOD@_ERR �wNJ�/�&PDUS_IZ  | ^���4>,5WRD� ?�E^� � guest|&l?~?�?�?�?�?�=DSCDMNGR�P 2x�E0�^| wd|&�KD	P01�.00 8C �  A  %�  

@�?@}�D�9 �������������hg@1g@�����XSM  �?G_�  �P�SO��ygG�E����R���{O��?@�@�D�0
�ZD�O�{g@��@U-w@�k@ew@��O+�+X�I0�+Sy*�d7OIO[OmO�;_GWROU�0y9@��2	�1.C�XQU�PD  Z5��T�PTY�`=�� TTP_AUT�H 1z; <�!iPenda�n�7Hn�/VP �!KAREL:�*HoQo|'nbK�Cxo�o^op`VI�SION SET �P�o�o�g�o'mc K9c]�������~dCTRL �{=&BD|!x �$�FFF�9E3�\FR�S:DEFAUL�TV�FANU�C Web Se/rvery*
Zd T?f4�|̏ޏ�����&��$WR_CON�FIG |�; �oV��!IDL_�CPU_PCu��|!B�_�� B;����MIN��D1� ?����GNR_IO1:2| 8���NPT_SIMW_DOΖ6��STAL_SCR�NΖ ��XINT�PMODNTOL8�؛��RTY�8ݖ�``ENB��R�|�OLNK 1};h0����į֯�������MAST�E͐�^��SLAV�E ~?;�RA?MCACHE*�"�}OaO_CFGl������UO`n���CMT_OPu�В:�³YCLk���o�_?ASG 1�7F1
 �1�C�U�g� yϋϝϯ���������p	����NUM9359
��IPi�{�RTRY_CNͿ�����Q93���5 �������J�\0���\0��P_MEMB?ERS 2��97Pk $������}���(逐RCA_�ACC 2��[�  QfNN �4� !c� _gp 6�zA.5B�o`v�%B  �_� 8�| /��� �3��X�BUF�001 2��[=� ��u3V�����u4u4�  ��u5u5���� u1u�1� �@u3u~P��`u:u:|!�tBtp�  � @~	� `u9u9��u7u7| �u8}u4A�u6u6| ��� u2u2Z_ 	�@y�`Y���q��y��u1�8�<Hp�	`�k�x�C�1h} �Hh�(��F!/`u1�0�DA�u2��_A�u3�T� X�u=�u=7P� i�N��@u o``a���	�`c�)�:���  u�3��u1�N{�u2p�3�hC �C91NNY�fU�  U����u0u�P������ y�@u1�a\н��3�h��0�8��sWu0�H�P�� ����2�������ns����#�5��G�Y�k�}�����XQ{��@�4����X����7 >���d(��?�`5���r�p���<����cм�@��Gn�/0HD�7I[m� y\�������3��( 22!HQ(-2a" 6-2AHSLOHRY HRa�loHRyHR Q"�d��d��d�� d��"��d���d��4�� �2:4���2
4���2�� �2��2*4!�b�4! �b! �b HQ0!5B4 /�@I"�@�4X#_@:4h#  p#w@y"� �  �B*4�!�B� �B��  
4�#� JD�#� �"�24��DX䊱2���]14�<�HQHP<�HP+T.QВX�HIuS�↲[ �v�� 2020-1'1-0�3{����_x�_�_wA $ ����_�_�_oo*o{�Q�g9hXt3yT9? %  ?.ouo �o�o�o�o�o�o�o�<bf�`h_zS��-�1PJ��-  M}�� # * {��6P(Qt�  1 �|0 : QtH�Qt��,R��5Q`Qth�QtpQtxQt�Qt��Qt�Qt�Qt�Qt��Qt�Qt��P��` )  EQAezd3y_x�Pp��EXr;^r7�|0C�� ��xp!  7�������~ , �p�+�.Q�Dd0G8-2�1�Hp_p���!�3�E��W�i�{�����P�4�؅5-2\31w6QQd��ϒHp;�bPp�ϒXp0.�Q�B6P4�
��!�3�E�W�i�B���v���B0x:��`Ԙ6`@[Pp��Z�Xp��a�  9 �|26P  " +xp9 ^��ߒ�� ߒl�ϒt�ˢ|�ˢ���8F�]������`(��ˢ�������!_��ˢ�p�^��;qK�pߒCY� R_d_�𬿾�п�Z)  Cۿ��*�<�N�<oNn*�p�ЊϜϮ��� ��������,�,|�1.�P��2 
 �SHp0:�OPr= �XrzЅ  ' %$|0;�� <��xp ��\��҉��� ��t� ��|��҄��Ҍ��Ҕ� �Ҝ��Ҥ��Ҭ��Ҵ�|���p,  G��
��E�p.\�������& #4��� W7 	|0Wp# U'k�Axp-ƀI�� ���������֘�X�p�N�p+�rՏ0����� R7�I�[� m������������Ǘ �Ԓ�Hp����XpT�҅ #�9��(``A��:L^p������6r��a�����9�Xp�҅ ��|0����;,��͠��͠����ҡ������ � \��͠��5������ ��p�W� �p CY � w��������Yt /'/9/K/]/o/]�o�9/�/�/�/ �/??%?7?I?7߶���c Q n�1s�3 �4(�40 �q Q8�4@�4H��4P�4X�4`�4h��4p�4x�4��4���4��4��4��4�z�4��4� r Qÿ`�#��A�W �4yB�0yB�0^�4�2 �0�2�0�2�0�2�0�2 �0�2�0�2�0�2�0�2 @�2
@�2@�2@�2 "@�2*@�22@�2:@�20��TO-wxC�xCY_ k_}_�_�_�_�_�_����z8U�4b�0b�0db�0V�49b4�T_ Yoko}o�o�o�o��*z8,�4-�4/�44� �0�"�0�"�0�"�0�""�0:�4ϑ�1>�4Er��0Er�0pr�0���0F��4��BJD}r@M*DO&DQ.DS6Db�h�I_CFG 2��� H
C�ycle Tim�e!Busy>'Idl�r�t�mi�2'��Up�v�qRe�ad�wDow������sCo�un�!	Num� �r�s�|+�� �Z�h�PROG�r툝��)/�softpart�/genlink�?current�=menupage,1133,�������/�
�"h�S�DT_ISOLCW  ��T�;���$J23_DS�P_ENB  �e����INC Q���#s�A�? ��=���<#�
<r�͙:�oi�u�` �$�+��OB���C�������E�G_�GROUP 1��e��< A���͑~)��3�?(��Я�!���/�@�S�e�w���'��=�G_IN_AU�T�pT�����POS�REM�_�KANJ?I_MASK�׺�KARELMONG ����"yN� g�yϋϝϯϲ�%²�%�����$��쿾��KCL_LǰN�U�p�$KEYLOGGING�0��������LAN�GUAGE ��m��DE?FAULT {ѰqLD�q������(F�����G�Ҏ���[��3 �� �� '�g  �[���>�L�;���
$�(UT1:\��D� F�S�e� w�������������(
FRA:\�RSCH2ﲾLN�_DISP �ట��㯹�OCT3OL��!Dz��n��ɑ��GBOOK ���d��������	-?�Qcs����	a	���ٍ�H��<�Ñ���_BUFF 2��e� �2 ���M�0�L^ ��������  /-/$/6/H/Z/�/~/�/�/���DCS #���ё[0	���sW��ݷC+��x��6B�뽔|��%?  A���>��A?���>
���� �IO 2��� !�p�?�p���?�? �?�?�?�?�?O$O4O FOXOlO|O�O�O�O�O��O�O�O__0_D_����ER_ITMb�d���_�_�_�_�_ �_	oo-o?oQocouo �o�o�o�o�o�o�o�k9tPSEVΰ��.nVTYPb��_mp�}�RST$���%SCRN_FLW 2�}=���� ��)�;�M�_�q���TP:�b�\r��NGNAM����m��$7UPS`�GI�p������_LOA�DJ�G %��%�J%qTUP	�R�A#�/���MAXU�ALRM!�б� �瞕
E��_PRD�а ��E�Cc����k7��k��P 2��� �Z$	���ΰ�ΰ#������$��!�Z� �H���t�������� ί��+�=� �a�L� ��h�z�����߿ʿ� ���9�$�]�@�Rϓ� ~ϷϢ���������� 5��*�k�Vߏ�z߳� �ߨ���������C� .�g�R������� ��������?�*�c� u�X������������� ��;M0q\��>�DBGDEF ��������� �_LDXDISA�ˀ���1E�EMO_{APŀE ?��
 ���0�BTfx��E�F�RQ_CFG �����A ��@i����<��d%��/��ؒ�����*T /V" **:_"��R/ d(����/�/�/�/�/ �/�/?5?���^?TP`O?�?s<�=�<,(3? �?���?O�?+OO<O aOHO�OlO�O�O�O�O��O__�O9_;�IS�C 1���E  � �?�_���_��_�_��_E_WR_MSTR� �-}eSCD 1���_fo�_ �ouo�o�o�o�o�o �o,P;t_� �������� :�%�7�p�[������ ��܏Ǐ����6�!� Z�E�~�i�������؟ ß��� ��D�/�T� z�e�����¯���ѯ 
����@�+�d�O��� s��������Ϳ���*��N�9�r�oMK���&m���$M�LTARM��:9'�� x3� ����į METPU�� R��.iND�SP_ADCOLx�� �CMNT1� $�FNM�Q�"�FSTLIr�c�` �&n�������|��$�POSCF��=\�PRPMP����ST/�1�&k 4�#�
a�v1a� q��]������� �������A�#�5�w� Y�k�����������$��SING_CHK�  u�$MODA��_[�˯��DEV 	�
	�MC:QHSI�ZE�P�TA�SK %�
%$�12345678�9 ��TRI�G 1�&k l ��~9M~=��YP�~53E�M_INF 1��9+`)AT?&FV0E0R��)�E0V1&�A3&B1&D2�&S0&C1S0}=�)ATZ�/$H!/I/�=q/ (Ay/�/\/�/�/�/�/ � ?���	/ z?-/�?�/�?�?�/�? �?O.OORO??�O ;?M?_?�O�?�?_=O *_�O�?`__�_k_�_ �_mO�_�O�O�O�O8o �O\o�_mo�oE_�oqo �o�o�o�_�_F�_ oo��So��o� ��o��B�)�f�x� +��Oas���� �,�c�P��t�/���𪟑�ΟJNITO�R��G ?e  � 	EXEC�1i��2�3�4��5�� �7�8
�9i����|�� |�"�|�.�|�:�|�F� |�R�|�^�|�j�|�v��|�2��2��2��2���2��2��2˨2�ר2�2�3��3�3"�R_GRP_SV 1��� (m���	����jv�
�e���&|��x�Ͼ���L�_D�m��׳ION_D�B' �+c�  K�c��@��%���c�h@ĐN ���J%�)���-u�d1: RSCH�\ݟ�ϰ�"�PL_NAME !�����!R-2�000iC/12�5L, Hand�lingTools  \�#�RR2��� 1��(��@��R� d��'�9�K�]�o߁� �ߥ߷���������� #�5�G�Y�k�}���<2#���������@&�8�J�\�n�<<�� �������������(:L^��|� � �� � ��  ��  A�  B� UT� ���
� �� ~���  ��� �� B� z� $�C���C��P E�;� E@ D�����D� ��8� ���  ��F
E�)>g+�E(� :9Z��H�%Z!fn/ W}��Y"JJ � =����>�>�+��(#�P0'%��(/2!&!F! b%J!%2%F%F!&!%Pf6)�%J!m� N+ 2%J!&�!�J2(��$I"�,1&S�)?�$?0'� �� a2��h?n1b1F%n?�3F!��� f&!�=�g�a �3�1f?�3�`�3|�?�6Fp E"0B�?�3�4F�?}6�>BO|7�bO�N� �E$E��L�E������� C � �O�K��d�C �D�O Y�O"_0W�@��8B]S��W%n__�_KV �X�_�Z�Ap� ��S������_�_	o�W��P��TB�i���Wogl���U	`�_�o�o|�o}a:�oA���o�o~;`\�)r �=f�_O:w|�l~{ �_�X�����t���R�� 1����R��bl6� Ē��� @�%?� v����?��v���@��6�Z1v�)�;��	l��	 � ~�� �,�^��|������ � s � � �䂱�K�l�,K���K���2KI+�KG0�K �U�����O=���@6@� t�@�X@�I�b�������N����
���ՙ�����_�����v�1a��k�ô� "����  �X�ￒ{4������r� ��  �����bW|2��>�T��f������	'� �� ��I� ��  ��Q�:��ÈƯÈ=��9�ޥ*�@��� �`��*�`�e4�8�[�p�  't���<S���?��b����^���C��B� C�4� ��B"ʱ��N��}�α����%���B�P� *u�m&p�F���kπ	���zϳϞϰ����5~ ������� �,0�:�d  >��?�ffA_$�6��� w`k�}�+��80��ߡ�?�R�$����(0���P����@�΃΄8�����Qa�;�x5;��0�;�i;�du�;�t�<!���C�R߄�`���&p�?fff?�?&���Nd@��A{#��@�o[�� 0��{���v���t� ��d纄U�*��N�9� r�]�������������0���F.p��,���P��q��C�?E&tPC�3�1�3̓ ��<'`K ]���`��� ��g-/�T/�x/�/ �/�/M��/�/o/?�/�,??P?;?�aA�x4�P�R�?AJ?�?F8xA�/C<?���?��?OO0������W0OC�T��` #Ca-O*�4��0�1��Ab�ܮ���bC�@_;CLn�B�A�Q�>�V�.È�����Y�\���
}OOc��Q���hQ�@�G��B=�
?h����O/`��W����ɰ�B/�
=�������=2MK�=�J�6XLI�H��Y
H}��A��12ML�j�LLPBh�H:��HK��n_�P	bL ��2J��H���H+UZBu2O�__�_	o�_-o oQo<ouo`o�o�o�o �o�o�o�o;& 8q\����� ����7�"�[�F� �j�������ُď�� �!��E�0�U�{�f� ����ß���ҟ��� �A�,�e�P���t���������ί��G�y��� C�a�?>;� Ĉ��]�d�OCVF酿���I[<Կ�@��Kտؿ� 
E�� �ƿK�z�@(�A�_�hM�����~����N���nπϪ�3lC�8�ϬϺ¢�������t�.3��}����k���q'�3�JJ��^�@L߂�pߦߔ��5P>�	P�����T��07�"�[�F��a�h����{������  fU���%��I� 4�m�����������������
��)�Z,  ( 5�{0HB�~�����  2 �E�G!�3E�L�n��q�5B��0�w1Q�C�l@�1  @Q�L�0 k}Џb��6��}Ӥ���//�//?�@#�8�4�y�0e��4�;
 0/�/�/�/�/�/�/ �/?#?5?G?Y?k?}?��J�2����V{H���$MR_CA�BLE 2���_ ���T��@P@PA? PA�1~�1�  ´ ��0C�06!O4>��B����rS�� ��6!K�p(� �����?�6��,  �� (� l6#N�/HB����)x� t� BR�eO�BZx,O>L<N@�` �L�D�߶B�%lhB�J�� . BC�͸�]�E�?�3 �O���O��O�O__  _�_�_V_�_z_�_�_ �_�_�_�_o
oo�o�|oRo�o�dE��  B��t�o��o
q�B����y�a�� ������`��� �ՠ���@��������7p��;p�?p� ����@�������7p�Kp�Op���3083/11|�l�3OM ��9����K i� �Z%% �2345678901��u ���qR6 �6 ;6 6!�
�w�mno�t sent *�K�6!�W���TESTFECS�ALGR  egD�;d��a!�
��� ��ЭD�3�l���ŏ׏� 9UD�1:\maint�enances.�xmYD,��kp*��DEFAUL�T��2GRP 2���z  p  ����d6& � �%!1st �cleaning� of cont�. vG�ilat�ion 56��Bԓ�@ޑ��+�a���"�4�F��m��G�w� %��me�ch��cal c�heckW�  ����C �������֯����[�w��o���roller�������ů�����п�1�Bas�ic quarterlyD�W�i��,��V�h�zόϞ�)�cMw���6 "8��!6 �����M�"��4�F�Xߧ�6!%C ;����ϸ���������
��k�}�Gr�ease bal~�r bush+���}���ߪ����h��/�A�C��geu��.L�t�y��  	3d�2� :�A��	��n���������}��
�gG��6&f�B��-6 ���]�@2DVhz}�
��cabl��6"�� ��@���
!� ,>�������������/}�Overh�au�ϕ�@B  !x�J!Q/���~/ �/�/�/�/�$o/�/�h�o? m/B?T?f? x?�?�/�?�/?!?�? OO,O>OPO�?tO�? �?�?�O�O�O�O_SO �O:_�O)_�O�_�_�_ �_�__�_ oO_$os_ HoZolo~o�o�_�oo o�o9o 2DV �oz�o�o��o�� �
��k@���v� �������Џ�1�� U�g�<���`�r����� ����̟�-��Q�&� 8�J�\�n������� �������"�4��� X�����˯����Ŀֿ �7����m�ϑ�f� xϊϜϮ�������3� �W�,�>�P�b�t��� ������������� (�:��^�߿ߔ��� �������� �O�$�s� ��Z���~��������� ���9�K� o�DV hz������� 5
.@R�v �������/8/�\	 T/I/ [/m/��/��+�-�/ �/�/�/�/�/<??? V?H?�?x?j?|?�?�? �?�?�?8OOORODO �OtOfOxO�O�O�O�O�\ ̼?� ; @\ z/Q_ c_u_\=_�_�_�_\w*�_** Q V�P�Oo,o>o obo8to�o�o���� �_�o�o�o�o1C U�o�o�o)��� �	��-�w�� u������m�Ϗ�� =�O�a���M�_�q�3�@��������\\��$MR_HIS�T 2�U��� 
 \d$ 2�34567890�1$�,���R#�9 ]����L�~�[ݯ� ���ʯ7�I�[��$� r�����l�ٿ����� ƿ3��W�i� ύ�D� ����z��Ϟ����� A���e�w�.ߛ�Q� ��SKCFMAP � U���R��Q��߳�ONREL  ���������EXC/FENB��
�Ӳ���FNC��JO�GOVLIM��d��g��KEY��zj�s�_PAN�ظ����RUNZ����SFSPDTY�P>�	��SIGN|���T1MOT\�����_CE_G�RP 1�U ���4 �_h�Q�U��� ������x������� ��?��4u,�� b����)� "_��|�p����/��PD�_THRSHD { Q�F@ )�QZ_EDIT�������TCOM_C_FG 1���!�؏/�/�/ 
p!_A�RC_���I�T�_MN_MODE����)�UAP_�CPL�/-�NOCHECK ?��/ �� M?_? q?�?�?�?�?�?�?�?�OO%O7OIO[O��N�O_WAIT_L���e'/�ODRDS�P�#��)�OFFS?ET_CAR[ �/��FDIS�O�CS_�A� ARK��f)O�PEN_FILE��@��!f&� OPT?ION_IO{���QPM_PRG �%��%$�_�_-SWmOP�?��ч  ���U���� ; �Ј �Q��P9'�Q	 �Q��Q�Q�zD��@RG�_DSBL  �����No��OR?IENTTO��?"�C�����A �BUT_SIM_DYW������@V�@L�CT �����*Q��$dQ�Z�dQ�<�b�c_PEX� �On�dRAT�' d)���d�@UP ��m�!ݐ�QcI���y�$PARA�M28��(��@�c �`/����%�7� I�[�m��������Ǐ ُ����!�3�E�Q�2�t���������Ο �����Q�<c�@� R�d�v���������Я@����������O���  ��  ���  A�  �BC�[ B�{s���3�H7��  �Y�?�>�BC�zC���z`yaQ�P �E;� EE D�	���M�Dn�����n������  �������E���Ѳ�gӳEc(�ȳ��Z��@Z�Ͷ�ɲ��/�� %�2�B��ʱ��b�Ȳ�>̅Ζ{���m�Ӱ���ÎP���ū���������
� ���������������(��2���m��NӰ�� ��ε^т���ȕ�������Bٮ�̳����ǂ�}���	��Ȁ��
����<����Ѓ����:���� 0l�n��l��`��~�>h�Fp Eʰ�����v�F3�%�� ��$炱
�4�+�0�&AB�g�y��d#�����������J�J�-CW%P�@��`X4^T
Ap?��g����q[�� ��BZ��2 ��P�mB3	`�HBTf%:��o�a����3 B�`�Z��2�� Ia/&+(I/ /m//�j/�/�/�/�F�r�pO�7p1�!�(�!���t0l�6!dA`��� @��?>�"1�G�?m@"1xb�˴x�"�P>;�	l22�	�P *0� ��,^L0M0k0��� � s �� � ��2� H���9H�H���H`�H^yH�R�,�hW��?�<� C�PB�C�ʰC4D;0O�#�9W�� ��k��}`�ʰ>A"O4O�FO�#�B<�{��KA��)O �"j��OK@���C�'$/2�?��? Q�V�/�0_�%	'� �� NRI� ��  ��MJ=����r_�[R@��_�P�N"a�_8["b�/�O�'N�`o  !'�`4d�1[@B:�B�}`
BoOAoSo -� O }�
A�8��`%�>�B�&B� �f ����Q�e���/��/;&_J\pOU�50`P�u�a�u E,KB:z�L2�1�D�?�ff�����t �)�[q8XK@?�M�?��.1Rz(K@{�P���y�1�z3z4�Sj����Zq;��x5;��0;��i;�du;�t�<!�ڲ?���04�S22�?offf?�P?&,��Wt@��A=#B�@�o[J�KI �b'���[p"5�� 7�� �f4�֟������ 	�B�-�f�x�c����� ��ү����m������4P��E C�۴r���?�����Ŀ��� ӿ���	�B�-�f�/ �ϕ�W�M?���7� � s�$�6�H�Z���o߁߀ߴߟ�����������A�$� �6�C���[���텹���?Ƀ؉�����KI�mرS�W��C� p�` Ca���ʣ����F�@I��Zn��bC@_;�CLn�BA�Q�>V���È����Y��\���
�)�����Q��h�Q�@�G�B=?�
?h�â�� ���W����ɰ�B/
=����Ɗ=JM�K�=�J6X�LI�H�Y
�H}��A�1�JML�jL�LPBhH:���HK�, 	�bL �2J���H��H+?UZBu�� ��|������ !1WB{f� ������// A/,/e/P/�/t/�/�/ �/�/�/?�/+??O? :?L?�?p?�?�?�?�? �?�?O'OOKO6OoO ZO�O~O�O�O�O�O�O _�O5_ _Y_D_i_�_8z_�_�YGϭ�_�_� C�a3��_ �爓�	ooCVF��1o8o����o�P���K�o�o� 
AE�o�oro�o�P(�Qϳ_�h�o����<*u�U�N��,��3lC�FXfr��r��t��.3��}��|k����q'�3�JJ�}�y
��.��(R�@�{�P�P�����ϭ� ���Ώ�����M�8�`��{]�l��q  fU ��H�џ���������`��L�:�p�^��v�0������ƫ)ZƯد  ( 5�'� ���<�*�`�N�����  2 E���ާ�E�L����ˍq��B�0�#��PC%��0��@�_���
��.�@�R�'������ϟϱ����ϧ�?)��ç��%���r}�v��
 �� ?�Q�c�u߇ߙ߽߫� ��������)��y����n{V{H���$PARAM_M�ENU ?�u��  �DEFPUL�S�l	WAIT�TMOUT��R�CV�� SH�ELL_WRK.�$CUR_STY�L�`��OPT����PTB����C���R_DECSN ��u� �B�T�f����� �������������,>gb�SSREL_ID  �u����vUSE_P�ROG %q�%8c�wCCR������y��_HOST7 !q�!���
T���9 �;u�_TIME���b�GDE�BUG� q�wGINP_FLMS�`̠�TR��PG�A� �|�+CyH��TYPEn�z�b\�/�/�/ �/�/?�/?"?K?F? X?j?�?�?�?�?�?�? �?�?#OO0OBOkOfO xO�O�O�O�O�O�O�O�__C_�WORD� ?	q�
 	�PR��cMA9I?��bSU�~ScTE\�c?X	���RCOL�e�Y�_@&�L�  �p��`���d�TRACE�CTL 1��u�{� |�o }p�� � ���|���:d	fDT �Q��u_`$`D� � u ���l`�pd�pac���b7a�aЂb0 ��bЂb	�rb��rb��pd�pd�pd�pdŪpd�pd�pd�pd�*pd�pd�pbE�cp �bp�bp�bp�bp��cE tpd̊pd�pd�pd��rbЪpd�pd�pd�pdԪpd�pd�pd�pd��pb\ !pb_ ��t�t߰�r�t��tpb^t^ *�t�t�t�t�u��t�t-��rs_�t_&t@t@t@TN�/s@6t@�d@*�tQ��s@�@ P�EP�P�� R�P���@�@�t@�t@��t@�t@�t@�t@�&�@.�@6�@ 
P�P�P�ӰR��sW@ "P�#P�$P�U%P�&P�'P�(P�)P�1P�2P���R�4P�5P�6P���R�UUP�VP�sP�tP�]u�g�tg�tUg&�g.�g6�g�Ug&�gn�gv�g~��g *�+蔟�g���g��g 7�8 �����&�ꒅ �ꒋ��F蔺�H
�I�J�Q ��P��M�g�h�i��j�k�l�m*�n�o�p�ŰR꒗�t/�\6�u>�Uutu&tu.tu6t)u�fGsuNv	pd��Uu�tu�u��u��Uu��u��u��u�Uu�u�tu�tu�tUu�tu�tu�tu&�Uu��u6�u�u&��u.�u>��suF�u�N�uV�u^�uf�u�n�u �pd�pd�*pd�pd�pd�pahb�C&tC�c� ��?�Ct�������� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� �����������'� 9�K�]�o��������� ��������#5G Yk}����� ��1CUg y������� 	//-/?/Q/c/u/�/ �/�/�(ha�%�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ���%�/>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r�������������&�8�J�\���$PGTRA�CELEN  �c�  ���b��x�_UP �����������x�_�CFG ���)��b������� ������ ��  ������DEFSP/D ����!� ��x�H_CON?FIG ç���g b��  dnMȇ� �!qP��b��x�IN~��TRL ������8�PES�]�����m\��x�LID������	�	LLB 1Ǿ]	 ��B&} B4M���!��f`��� <<7 �!?��� ������-// E/c/I/[/}/�/�/�/�/�*y???K?��D?�?t?�?�?�	G�RP 1�2�G�  ���
�b�A�PH���@B��A} D�	� Ap	@�r�$I4Imm �`�?�PN´�CiORKB�@�A�O{O�O��O�O�O�B��B�C5	_B_T^>_ <�oyQY_�_U_ �_�_�_�_�_q_�_4o �_DojoUo@z�c�ob�
o�ooo�o�o�o >)bM�q�������b:)�b�)
V7.1�0beta1� @�{@�?�A&�H�1=��C� CzB�O�D71� e�C�� b�ߛ� D�w�A@� �1B M@�1C6�1 �� �!�!#C�����B��0L ���%���0CRL���	����AK�33AFff@s�33BZ�z�!A��ffA�33@�����^�#E�N���b����O ��Fq���m������
�KNOW_M  ���SV �]
���oQ� c�u�Ɵ������ϯb��,MM�3�] ��M�	����C���:�����Ic�$@>� y�u�X��� MR�3��eT�J���b�C�c�U����OADB�ANFWD� S�T�11 1ϧ��?�4EOAT� with to�te�B@?�  ��L�33F����G�3F���fc�]�no8f�Ms� ���� �Iش��������� ��/�a�S�eߪ߉� ���߿�������L�c�<�2G��4/� � �<��X��03 n����<�4��������<�5�&�8�J��<�6g�y�����<�7 ��������<�8X1C<�MA'�-D�k��OVLD � c3��>�P�ARNUM  �J��\�39�SCH�	 �
IW5�iUPD�dE|���_CMP_���� K�6�'3��E�R_CHK����3�����RS8ư*��1_MO'�J(�_7/_�_RES_GF��c
���/d= �/�/�/�/???I? <?m?`?�?�?�?�?��#m��,�/�?�%�� �?OO�#�3OROWO �#f�rO�O�O�#��O �O�O�# �O__�#�_ /_N_S_�"V 1��J�/���P��`M"THR_IN�Rư��3�d�VM�ASS�_ Z�WM�N�_cMON_QUEUE �J�X3�[ � _�N��U!Nf:hQcENqDVat/piEXEo�pe�BE~``oQcO�PTIO]g}+T`P�ROGRAM %4j%S`�_8Rb?TASK_I��nOCFG �4ox�([pDATA��]�d{@�v2+ ���
���;�M� _�q��������ˏݏ^�zINFO��ը}(�ȓ�0�B�T�f�x� ��������ҟ���� �,�>�P�b�t�����4� �֨| �9Zq6PK_^q�dy �ۦENB� ꭮�
�i2�%�G^q2�� X,		!o=���q�����$U�!�����T֧�_EDIT ��d߿�WtWERF�L�h�S9�RGAD�J �κA�  <�?[ H��Q �Ta����K?�A�z���q<��~)%DIAG��`�Ϻ�	_¸�2�j���	HK`l���RBp>��UU@\x��*,�/.� **:7�'�9�Y���P>��� �@�u�ߴ��Yzu�8>��:�߀���߸��ߺQ�PA������g�%�7� �L�v�����������r����>���v����AP
�^� X�j������������� P��L60B�f ����(�$ �>�zt�  /�����l// h/R/L/^/�/�/�/�/ �/�/D?�/@?*?$?6? �?Z?�?�?�?�?O�? OO�?O�O2O�OnO hOzO�O�O�O�O�O�O�	w�_�o_�_�T�t$ �_�[�_�_�_o-oZ�PREF� �j���
~ �IORITY�g�ն�$�MPDSP0�a����gUTFvӾ�ODUCTCqeκ0o��OG���_TG�HrҺ�bHIBIT_DO��{TOENT 1��λ (!AF_INE�`epw!tcЉ�{�!ud��~!icm�]��bkXYc��μ���)� D�$�6����_�B�N���r��� �����̏	���-�?� &�c�J�����*�cc�	�j���%G_ݟ�yb�>�%�"�D�/N�˟@���������>�,  �``Ρ@���������e�0��Z0����#�5�����ENHANCE� 㺝��AЫd /���|��fId�Qocc��$�PORT_WNUM�c�e�$�_CARTR�E{�	�Z�SKS�TA�g2{SLGS6bp�	���Ù`�Unothin�g��zόϞ�7k>�T?EMP ��i���?Ub�_a_seibano� o� C�.�g�Rߋ�v߯ߚ� �߾���	���-��Q� <�u�`������� ������;�&�8�q� \��������������� ��7"[Fj���������VOERSI�`�g.� disab�le����SAVE� ��j	26�70H722��!������C 	��bA_+/�ce,/U/g/y/�/�*AD,��/˭K_p� 1�	�w ��:
W?+?�WB`URGET�Bp+~�qWFW0'q�d�j��fW^px4�a��W�RUP_DELA�Y ��k5R_?HOT %fV�a����?�5R_NORMAL�8�b�?<OGSEMIOAO�O@a_QSKIP�#���3x��O��O�O_ �M^]<_lS@_f_x_�_ P_�_�_�_�_�_�_�_ ,ooPoboto:o�o�o �o�o�o�o�o: L^$6���� �� ���6�H�Z�K3RA���Kh�H���t�_PARAMv�A2�K @g��@`�&j�2Cju��BÁC�&zձBt�BTIFy4��RCVTMOU�&���t�DC�R�#�I ���AE��ED�E܅vD���C��OB���(��Gţ����Љ�	����9�Ú�A�Ǖ�z�O��_ �;�x5;��0�;�i;�du�;�t�<!�� ذ���&���J� \�n���������ȯگ�������RDIO�_TYPE  ��-��ED��T_jx����X�BH�#�E��j����z� ��B����Ϻ� ������=�(�пn� mO��$_��������� ���4�"�X�Bׄω� �P߲ߠ��������� 
���T�v�{�ߜ� 6������������ >�`�e���6���2��� ��������:\� a��B���� � �$FK] ~������ � /BG/f(/z/h/ �/�/�/�/�/�/�/,/�R/C?�j�INT �2��9���4�G;� �?�;� ��?-�f�0 �?�;?O �/OO/OeOSO�OoO �O�O�O�O�O_�O�O =_+_a_O_�_�_}_�_ �_�_�_oo�_9o'o ]oKo�o�oyo�o�o�o �o�o�o5#Yf��EFPOS1 1��9�  x�AT HOME���Ճ��(�1���z��lu�
��Ż�ۿ�xߣ���(�={�5�}@N���=1?����?H�3�l���ABOVE �LEFT JAC�KP(�Ň��+^���H�~�Ff#����4��+�ɏ��|�~����ڍ@��<z���RIGH�����,^�@I���G��*;��"y��nʿ�ʏ܏��"�\� ��X�џl�������+���O��EO�pc�hange po�s�w�g��?���x=�̅��<<!H���%?�N�����n�MAf0 1���d��ɾI�/����E�<L�u'����C������ί�2���e���>g��࿊H�<ǘ����x4��!�"�8�F��3c���f��ʣ��
�ٿ5S�;j{��?3k���������At �Pallet S�top餡�o�����>�����=�9)D��?t8>[���(��6�H�a���p������վQ@����8xvտ�?T[��^��Ϡ�Ю���ٴ��q��d���>	�
�
E�e�bٿ��������&��8� 4|�r&���=�����6K�f���!�4�]zߐߞ�Ұ� 㡉s���6�9�Յg�����3�ⷿ�_a��!���'��p 6|�t��B��E=�Eȿ	��I������/���Fej��� ��<�M�8�q���� 0������������� 7��[mT� P�t��3 W�{�:�� p��/�A/�e/  /o/�/�/�/Z/�/~/ ?�/+?=?�/�/$?�?  ?�?D?�?h?�?O�? 'O�?KO�?oO
O�O�O @ORO�O�O�O_�O5_��O?_k_V_�_*U}u2 1�3_E__�_ �_!o'_Eo�_ioofo �o:o�o^o�o�o�o �o�oeP�$� H�l���+�� O��s�� �2�l�͏ ��񏌏���9�ԏ6� o�
���.���R�۟v� ����ԟ5� �Y���}� ���<���ׯr����� ���C�ޯ��<��� ����\�忀�	Ϥ�� ?�ڿc�����"ϫ�F� X�jϤ����)���M� ��q��nߧ�B���f� �ߊ��������m� X��,��P���t��� ���3���W���{�� (�:�t��������� ��A��>w�6 �Z�~���= (a�� �D� �z/�'/�K/� �
/D/�/�/�/d/�/ �/?�/?G?�/k??��?*?�?�_�T3 1��_`?r?�?*OONO T?rOO�O1O�O�OgO �O�O_�O8_�O�O�O 1_�_}_�_Q_�_u_�_ �_�_4o�_Xo�_|oo �o;oMo_o�o�o�o �oB�ofc�7 �[����� �b�M���!���E�Ώ i�ˏ���(�ÏL�� p���/�i�ʟ��� �����6�џ3�l�� ��+���O�دs����� ѯ2��V��z���� 9���Կo�����Ϸ� @�ۿ���9ϚυϾ� Y���}�ߡ��<��� `��τ�ߨ�C�U�g� �����&���J���n� 	�k��?���c���� ������	�j�U��� )���M���q����� 0��T��x%7 q�����> �;t�3�Wx��?�44 1��? ���W/B/{/��/ :/�/^/�/�/�/?�/ A?�/e? ??$?^?�? �?�?~?O�?+O�?(O aO�?�O O�ODO�OhO zO�O�O'__K_�Oo_ 
_�_._�_�_d_�_�_ o�_5o�_�_�_.o�o zo�oNo�oro�o�o�o 1�oU�oy�8 J\�����?� �c��`���4���X� �|������ď��_� J������B�˟f�ȟ ���%���I��m�� �,�f�ǯ��믆�� ��3�ί0�i����(� ��L�տp�����ο/� �S��w�ϛ�6Ϙ� ��l��ϐ�ߴ�=��� ����6ߗ߂߻�V��� z��� �9���]��� ����@�R�d���� ��#���G���k��h� ��<���`������A��*SYST�EM*��V9.1�0170 G9/�18/2019 A �  4���#51_T �  l $C�OMMENT �$ENABL�ED  $A�TPERCH�D�OUT_TYPEz� �INDX���	    	�TOL�HOM]E� Hi6q�w����� +i7q�p*<N �i8qq������`SMSKr�  $MAX�jEN�����i MOTE_CF�Gr T $d�$"" �#IO �*I, �!LOCA�L_OP�%�#ST�ART{!��i POwWERr m /FLAG� �"�"�r , �&$�DSB_SIGN�AL�"�"UP_C�ND�!�4�R�S232�% �� ��DEV�ICEUS�#SP�E �!PARIT�Y*4OPBITS��"FLOWCON�TRH �!TIME� �"CU�0M�"A�UXTASK�"INTERFACi4/TATU�0u � �SCHr 	 t��OLD_o0C_�SW"FREEF?ROMSIZ "� GET_DIR��	$UPDT_M�AP "� Td EN�B"EXP0JC!�`0FAUL@EV�!�RV_DAT�A�1
  $zd@E�1   ? �VALUyA> `FG?RP_ �"dA�  2
 �S�C�"	� �$�ITP_vB o$NUM�@OU�!~�CTOT_AX�1��CDSP�FJOG�LI�3FINE_sPCZ1�1OND�E�o!�@�6K+@_M�IR�ATP� TN�5XAPI 0!RE_EXXP2D�A5 .Q�"��APGmVBRKH��11FNC�@I:!C  �R#�R�BP!@�D�!�C1PBSOC��F� N�UDUMM�Y163�BSV_�CODE�!*3FS?PD_OVR |@��LDb	SOR$g N fF�P2g��@OV�ESFJjR3UNMc!!SFff�!�SUFRA|jTO~�4LCHDLYWRECOVd �@�WS @�P�e�@RO�3�QP_f`  � @� Su@NV�E� !OFS�`C�@ "FWD.a�d*a��Q�QU�PTR)1�o!_VQFDOQVMOB_CM�!<pB�@�BL_c S^rdq2ncV�1 "@s@�CFbG_wrXAMpSRp�0��u�b�_Mvp�2Mx�@�"�`T$CA�@��pD�R�pHBKX!A0F�IO%��!"�PPA	�5���E�-��u�"�bDVC_DBG #w�1A2w��b�!��1���s��y3���`ATIO� �1�0aU #�@�&CAB P" "P�d�1 �x!!�@_�00FS�UBCPU2PS�IN_0Hs�t"@1�D�ws�t�"�Q$HW_Cq �0S�$�|��wq
 @|@�$U�NIT�T����A�TTRI3@��PC�YCL#NECA�ۂBSFLTR_2_FI-#/9�"6!!{LP[CHK_�0�SCT4SF_��F1_��.���FS!1�r��CHA=��o�r�2n�RSD�`2�Q�;C1� _T�xPR�Oǀ6s�0EM _D�@�ST\�S�|@\��wp�DIAG1ER�AILAC��*�MF�@LO�P!�V4�BPS�B" #���skPRx�S$@ ��M�Cj�\0	�cFU�NC�R�1RINS_T$A ��m��1#RA~��@; �p��8p �t��WARBP�?CBLCUR��ǴaA����ø��DA�P0���ǳ��LD@�P�"�)��A��.�)�T�I:�IſA|@$C�E_RIA�1+2AF:�P91t��`zŋT2�C/C��qqOyI��9vDF_Ly �~bA�0LM�sFA>�`HRDYOBQ�`RG.�H��4Q 	�>��MULSE��3C�I��P��$JjJ�,bAg<kFAN_A�LMLV)3H�WR=NO�HARD !F�P�2��2Gф1�A��U_�`0FAU�0R�a��2TO_SBR �%���@�ڛ�l�u���_MPINF�`��������REG&NQV@��VD� NHtsFL}��R$Mʰ ��3I��p|@V�]�CMj�NFƑ !4��?pprk $�-!$Y��A��B�As � ��eSEG���C�P��AR�@�#�U2�S����rUAXE�GROBn�JRED�FWR�`2�Q_#��SSY�P��t�PE�SO�WRI�`��{�ST0�C�0�P
 `E��? ��)���"�@B���a��5��p�OTO�? �`ARY�C���˄="�0�FI{P�3$LI�NK��GTH���8@T_���a��6��BXYZ!B
7N-OFF�`��J��B�@b�r0�a)0@sFIʐ���0*3�Tb��D_J Z1|Bb��"��Х����8�Bg0�����CL�!bUDU	r��9*�TURJ�XP�4��b��X^��p�FL ��`����R6��30��Bq 1? K PM0D�U3S�-�I�8:�I�	CORQ���A ���wq-�xPOA�z!�b�$3C�A�$OV	E!��M�0!��8% ��8%��7&�16'$A6'@5$ANs���8!z� ��!/Pw ��!0%!�<'�%���%\#�AERQ��	.�E�`d@:��$A�!|@�����0�����AX�c|B �������Y5�e9� e9)�d:��d:, d:K  d:� d:+d:1�d6 ��a9��q9���9���9 ���9���9���9���9����9�1�9DEBUs�$n�z�⢢Ar�AB��.a#V�pr� 
�B���� �Ewq�G�Q�G)��G�� �G,�GK�G��G+��� z���sLAB��o�|�GROh���s��pB_ȡ �&{�'c� �КV�Q�8�U���VAND�.�@�$��!��g �q�{��'h��6h� NqTZмcY`VELΡ�$ca�kf�SERsVEY`�� $��ښ�A�!�`PO �bs�Ap��a �b�!���  $.�bTRQ��
�c.��`�gz�2�fX��?_  lX��qN�ERR�q�I�p8g`�$,qTOQ�$� AL�c4k�?v��G�e�%� �cRE>
�  ,�a�e��`�"RA�q 2g d�r-��|tn�` ��$, �͢��S2 ��aOC|���p  {�COUNT�� �_S�SFZN_wCFG�a 4x���T�p���Cs��@�vr �`��� ��@M=�!Ҡ�Հ0�#5!=�u�FAg��%u�y�X�u�Uq��$�d��P���`�HEL7��� 5� B_BA�S�RSR�V�"�S��B��1hw�U2*�3*�4*�5*��6*�7*�8hw��R�OO�op�� NL���AB�c ��A[CK�FIN�pT!��M�U����a���_P�Ut��OU�cP�~���ivb�}�?6T�PFWD_KAR�1q#� pRE�d��P8���s�QUE麠  ltЇ�IK��C�� �h`�SE�M�A���A��Aq�S�TYɔSO����D�IՑ{�7�u�>7��_�TM/�MANRQ�� END��$�KEYSWITCaH�-��~�HE�BEATM`�PE���LE0r�Q�P^�U�,�F��-�S�DO/_HOMx�Opѽ�EF� PRx9�0�|�֕Cx�O��p�q�OV_M�s�Y�IGOCM���A�bv�HK�� D$�G�Urs�M��G��X FORC �WcAR��yr�OM��  @�D���U��P��1z�]�|��3z�4�����US�pO=�L`��r��UNLO�t���ED�� �q�PHwDDN�a �`�BLOB  ^��SNPX_AS�� 0D�ADD|G�`�$SIZuq�$VA�PjuMU/LTIP�����A`� � A$�Ь�� ��S7��QC,py�FRIF����pS]�oɰ�i�N=F	�ODBU^�8`�zսӸ٥fw� �IA`N�������S�>�� � #�Ir�TEm��SGL1�T��^&)�J�S<G�2�STMTkc�P��o�BW 3�S�HOWk���BANw�TPU �+��h���pV� _GY�;  � $PC�P�p��#U1FB\�P��S�P��AԐ���VD���X�!� �qA00d1��9�@��9���9���9�57�U67�77�87�97�A7�B7�n�9�mQ:���9�F7��0��C��Р��]����w�1��1���1��1��1��1���1��1��1��1���26�2C�2P�2�]�2j�2w�2��2���2��2��2��2���2��2��2��2
��36�3C���]�U3j�3w�3��3��U3��3��3��3��U3��3��3��3��U46�4C�4P�4]�U4j�4w�4��4��U4��4��4��4��U4��4��4��4��U56�5C�5P�5]�U5j�5w�5��5��U5��5��5��5��U5��5��5��5��U66�6C�6P�6]�U6j�6w�6��6��U6��6��6��6��U6��6��6��6��U76�7C�7P�7=IU7JI7WI7dI7qIU7��7��7��7��U7��7��7��7����VP\�U�b"��¶P�
�Ҏa#� x $TOR f������r�`R�`ڀ�TQ_�pR�`Au�a�8�ndSmC��e�5f_U��@a�YS�Lfp�`$ �  #���$���ג�� ��<ld��VALU$�ߐ�2�a�hF]aID_YL���eHI�jIN�?$FILE_��d�#�$��CYeSA��q% h�P$pE_BLCK`�1rL�>:xD_CPUJy$�@Jy�/��otU�Y1�� �R & � �PW�p���ЫqLAq�S�p�t�q�tRUN_FLG�u �t�q�t0��u�q�t�q��uH ��t��t��T�22�_LI`�' w ��G_O��}:�P_EDI��f��T2��:�(B���ɲ�EqkР�`�BC=2#�) �(�$�0�p����:�FT����.ãTDC�pA��Q��ɀM�PÆفTHD�Ѐ���S��R��<���ERVE����ã�ፂ� �*X -$H�L�EN��U�ãH��R1A\���\`W_awsi1H��d2��MOBq��S��ҐI�1b�a0���TH�̛DEܕ���LACE�cCC8��1bp�_MA	�ۖ8���TCV�=��T�>�]�S��ړP�ၥ���JΠA��M����J��!�ڕǡ�T�2�������ٓ��JK�VK@\�� �����J��l�	�JJ�JJ�AAL	�?��?�9�d�=�5��p�N1d�Pp�/��dL��__��������CF�+ =`�PGROU�`Mᔹ���N��Ca���R�EQUIR�ƠE�BUx�D���$Tܐ2*�E�붎��Δ�, \B`t�AP�PR��CLb
$:K�N>�CLO��NɑS�c�ڕ
��L�- ���M׀�o���N��_MG�Ѩ�C#��%p�ȧ����BRK���NOLD�ƒ�R�TMO9����͢�J9���PA����������]���f���6.�7�.�?�@���.�# ��o�\��� ���PATH�ױѧ� ��t��ӎ��-3a���SCAx���?§�I�NG�UC�����C��UM�Y��p ����a#�2��2�H�~2�PAYLOA���J2L�PR_ANρs�L�p}�y�m�����R_F2LSHR���LO~�U�������ACRL_@����� �e�g�H�`�b$H��%�FL�EXA���J��/ P+£����.������JG�0 : T�f�됷���i�h��r�����F1��0�����ɟ۟���`E 	��-�?�Q�c�u��� ��7T�����D f ��̯ޯ���T�5X=a������% ���,�>�B�K�9��]�f�x�������1 �����ο�퀺PcATI󱥠EL� ���3��J�0�J�E��CTR �DT�N�Q6�HAND_VBbA�`��72 $�F2���m�cSWrC_�����3� $$M �����P���8���<� �5��6A�`j���aDI��A�̖`��A��AA��@��cp��D�˕D��P��G�p�IS�T�ǼA�ɼAN��DY�p<����4&E��I� �������l�������P6�?�H�Q�Z��c�l�uҩ�J��41 �0���� q�U<p��QASYM��@`	����3"a������_�����	�d�8 )�;�M�_�q�Jx�)����c�i��V_VI�r3�hp��`V_UANY��`s.#��J�� %rSU%r��)t��6tZv ����)�
���u�a2�:�2��HR���w�5�2�qT�N�D	I���O�t�2�p���6 > -BIaA -���'�J 5c5�M '0��0� �p 7 �[ �1ME�� hP��r7aT�pPT�` � ��x����$S�o`�}�����T�`�� �$DUMMY1�H�$PS_G RYF	 ��$ӆ��7FLA��YP�����$GLB_T �0�u�x�\��� H1�T�8 X+�뷂�SuT���SBR���M21_V��T$_SV_ER��Ob`LN�f�CL"�N�A� �O*��pGL�`EWβ�9 4����$Y"Z"W��頲�r�3AQ��VRD��]U��: �Nːޓ`$GIX0}$�� ����ʐ���; L���ab}$�FabE��NEARʙ NNF;�� TA�NCN���JsOG��� <� $JOINT�x� L���MSET��=  �E!�K� �S�"���� ��>�� E U�?���LOCK_FOx��1�pBGLVK3�GL�TEST_sXMA���EMPw����	� �Р$U�� 2:�ʓ/��;���0ՠ/�9P�C�E����P� $KA�R�M�sTPDRqA��m�d�VEC��~�h�IU/�<4�H=EנTOOL���VRE��IS3��ò6Q�D ACH���=��O�Ѐ��3>!��SI1� � @$RAIL__BOXE�s�oROBO �?�s�?HOWWAR-��<Ѐ�ROLMۂEŀ�!�V��!�8 ��O�_F� !s�HT'ML5�q �%���tݱ��?p�
�R��O��@�� y�}���v��OU��A d���+�97a!2�!Р$PIP�N�����ݱV /�����COR�DEDՠ�п�8�XIT��)�p� O7� B D �OBSA%3ՠ^�MѼ�p�M�a`'1SYSM��ADR&1�px�TC}H�0 C ,�SEN�r]�Aܡ_���Դ!AՒVWV�AS�D � �s����uPREV_�RT`Q$EDI}T��VSHWR�!�:������`D�b���5�.!$H�EADra�pO��a��KE����CPS�PDf�JMPj�Ld�u@�R� �EU�TR��I
�S&2Cl0�NE��'1b7TIC)K�aM[�����{HN0�F @W�8��%n�_GP����^�STY���LO�"�� ������G �t 
��G��%$����=:�S !�$q g��$��P�P��SQUg���aTERC|�!G�=S�$H �F�@�'��'g��(0O}��p�R IZ����ρPR3�܁����sPUq+_DO@�ֹ�XS��K�vAXiIJ i�4�UR� ��'2&���x֗1� _,����ET�Pޢf�J�UI�F�WJ�A�A�QÄ9�>0 ����SR4Il ���9��:�6�2 GIILAG LQGLaF^x�I^H��R|C��C�`Zolo~o�d��SC
�� J hs�DS���SP!�x%A	TO@�2,��⿂�ADDRES��B�
�SHIF�#&�_W2CH&0t�I)���!�TU)�I�1 �K��CUSTOT�5�V��I�L��P�!�P
	�
a"qV��;U�M \������I�<���W2C��C��):��l�W1�TXSCREEO��N�pe�TINA�����4��ь�"�PO T��i��� h�E��6X��X�4�RRO*PU���`��1�F���UE��P ���P���S����RS	M��NU<е��vaA�pS_ē�FcqA�I��Gc�Cʢ]B�4 �2O�0UE�TQp�y��F GMTmp%LGqgU�Oz���/BBL_�W��U��R �I�!RO��-RLE�"8S%��"7T�RIGHASBRD<{��!CKGR��iU�T=�hWeQWIDT�H�+�E� �큭�oD�UIx�EY� �T�S��D�-��BACK+�ۂ�U��[�FO*��WL[AB6?([�I�΢$UR+�`?A�I_a�HA T 8�qU�_N��"?bb�R��Т��ˁa�R,aO�!U�U�����bPUMP�cRޢP�L�UM�co� ERVH���еPP?��TVY�� GE b&�� C�&W�LP�e�E��=!)�g\�
x]!
xװ	yU5{6{7{8�b���p� ?�k4��ױ�ȡS��U�QUS=R��W <��a�1U��#�FO� �PRI�m��{q�p�TRIP	�m��UNDO�X�`n��pP7�O)�&�� �� Y:b�pG V�Ti�+!�!&5�OS��J�R� B!���1�Z������q�H��a'�U�a1�[z�����C�b�!�OFFT��2�\6���O �� 1Zs���[s�GU��P�{�-�8(!7��QSUB�N�@SRTs��]��T�u���OR�}�RAU� ~�T����c�9_�Е�^ |���OWN$���$S#RC(@�@l�D����MPFI$�S!� ESP'���0���c�<�gɲ �����A_� `ÀWO2������COṔ$� &�_���w���~�WA
�C���[�1��Z�ɲ�0��C�1 �`�2SHADOW�l ��͡_UNSC�A��ͣ�TڣDGD<�e�EGACq�75H�G�2a:bh'STE4Q:�Ox`�d��PE�bgVW:���TRG� �A�b ���0�MOVqE(C��ANG�D���؃������LIM_X̃��҃����ı����CK��p� ����VqFi ~�`�VCCM�j��c�2C^�RAO�p@�z�� 5�NFA�i���E�a�p�G� APb��&�D�E^�1�.E��Ad�� ��z� Dű͎�dcpC���GDRI����j�V������� D�tMY_UBY�tE�q�z�)A����0<�@ر�O�P�_�$�a�L1BMv4Q$��DEY��cEXP5C��MU��1X7���v@USkAv �p_R�1���p� ��=G�PACI�g� 󑋴��؃�җ��ҩC���RETb�!q�:�8���ҙ�e � i�EGk�P�29���Ra����f�P�`A�Q]�	4v�HR6�SW��Ò<��� O�q�QA(� ��EzpU<�]�n<�$C��HKA�g�`�ꏱ� ���0��EAN��Z�A`�弯���MRCV�Ah� ��`O5�MA`C3	=��6�=�REFW_�F�1񵲸�� �pB���S���d���F���_������4��4D2Ҟ0Z�9��Di �H�l0z�#�q�?$GROUv ���0�mE�w�dO�,!2�e�@�0m08�Pf`�#,!�R@� UL��eg6�CаUah��� NT1�����na��q�� LK�
[�P
na�q1�T�nDDj tÀMDi�AP_HUZ���V�SA��CMP(@FP\um]_t!RĐS!��X�Z���VGF����k�� �`M�pAP0�U�F_&@v�/��uROKP�2�7դ`F��P���URE�RA&��R	I��_I� g���������ȹ�҃�IN"��HT$#ȜPV��ײ?��#{S�%W��'熡`�Á���-9��LO������#P9�\1uqNS=I�VIA_Z��0�l �+PHDR =�P$JOupR��$Z_UP|԰-BZ_LOW�5�y1�GaRӰ[AL P��W�B��1y1- \@Ĺg�0Ax0���m�� 0�PA�Q= �CACHc4P1�(EO1��DI�a���CJӱI�F�1pET<P�oF'$HOA`*� -@��öb"�FP�R`����aT�VP3�<]��B_SIZZ��D�Zg��H�1�G��|SM�PZg�IMG[��N0ADMYw�MRE�SmRWGPM��N�D����ASYNB{UF��VRTD�U��TQ�COLE_2�D״�U2܀C�U��[@Q���UECCU&�VEM�(EbnGVIRCMQ�U�S�b�Q&0LA+���(���<�AG�YR��X#YZ� ����Wj�h��!~dS�,`TE���I�Mea�VGb�cEGRWABBn�Y7� E�>n����CKL�AS*@��AK@o�  �`T4��@Ģ�*�$As��p A�v!��0b�#LuT� ����7��r#�Ist'��Kf��BG_LEVE����PK��Mf�6PGI<pNO7��ћNT7rHO���q � w�_� �Pb�vS�0���RO��ACCE��]�#�VR_c��M`$�����6�pARE�PA��S��� Dq�REM_B��d �b_JMP�  ��rt�$S!S��t�0GzQ@'s ��[ASoPJ6}Nڅ�VLEX=v�tȢ����� �DDR��$��Ӡ�}��\���P2Fu'� i!?�V_�MV_PI�Su�T ��z���j ��F�0�Z������y��!���!̪�h�GAɕ��LO9O~���JCB��~w��C���@֣PLANҲqB�r�F"SO���P\�MQ�)�Ń���S+К�P����!P�@nB�!��PâT?���PRKE�N�VAsNC�?R_O�@v (B���ɳ�Sp��S�rR_A�� w 4R�!��ΰ�p��k�x h��ࢉ}1�W�OFF�v�F\`eDEA�j�
�P�PSKsDM8���� w ���@|'�ry < ��-��UMMYj2�D2��_��CUS��U��z� $� TIT��$PR�+�OPLG�t3SFD�\�{p����P&�SMEO�|Ђ�K�J;�����0Q_�E�}�ЂX���0��@��XS�~ x�0M�SPD_���1�`P��`�S40NB�2LNTK3�M�>4�p�C�0#���1Ҷ�'n$�XVR��b�X�T6�
�ZABC=�K��-z~�
s��ZIP���Ђ�pLV�CL�w�~���ZMPCF�Ղ~���3�V�?DMY_LNϰı�D��� �ԃ �$�A ��CMC�M^ C�CCART�_G��P8� '$Je�_�D�Ak� |�u� �� _�R�Y��z��UX�a
�UXEUL��ap���������������d�FT�F�k�%�m�����G� ��w�?�Y�0�D�` � 8 �$R[PU2��EgIGH�X�?(� �����c�>� �0�pf�q!��$B� �0<}2SHIF����RV=�F����	$��6�C�0`�U�f��0�
Ks&�D&6TRb �V�Q���kPHB�K� ,�� z�������0F�� 5 1 �����  x�I ���	 ���  ��gR� &�J�n�	/� -/�Q/�u/�/"/4/ n/�/�/�/�/?�/;? �/8?q??�?0?�?T? �?�?�?�?�?7O"O[O �?OO�O>O�O�OtO �O�O!_�OE_W_�O_ >_�_�_�_^_�_�_o �_oAo�_eo o�o$o �o�oZolo�o�o+ �oO�osp�D �h���'��� �o�Z���.���R�ۏ v�؏���5�ЏY�� }���*�<�v�ן�� �����C�ޟ@�y�� ��8���\�������� ޯ?�*�c�����"��� F����|�Ϡ�)�Ŀ M�_����Fϧϒ��� f��ϊ�߮��I��� m�ߑ�,ߵ���b�t� �����3���W���{���x���6 1�S�e����A� G�e� ���$�����Z� ��~���+������ $�p�D�h� ��'�K�o
 �.@R���/ �5/�Y/�V/�/*/ �/N/�/r/�/�/�/�/ �/U?@?y??�?8?�? \?�?�?�?O�??O�? cO�?O"O\O�O�O�O |O_�O)_�O&___�O �__�_B_�_f_x_�_ �_%ooIo�_moo�o ,o�o�obo�o�o�o 3�o�o�o,�x� L�p���/�� S��w����6�H�Z� ���������=�؏a� ��^���2���V�ߟz� �������]�H��� ���@�ɯd�Ư���� #���G��k���*� d�ſ��鿄�Ϩ�1� ̿.�g�ϋ�&ϯ�J�x�Ϲ���7 1�� �ϒ���J�5�n�tϒ� -߶�Q߳��߇��� 4���X�����Q�� ����q�������� T���x����7���[� m����>��b ���!��W�{ �(���!� m�A�e��� $/�H/�l//�/+/ =/O/�/�/�/?�/2? �/V?�/S?�?'?�?K? �?o?�?�?�?�?�?RO =OvOO�O5O�OYO�O �O�O_�O<_�O`_�O __Y_�_�_�_y_o �_&o�_#o\o�_�oo �o?o�ocouo�o�o" F�oj�)� �_����0�� ��)���u���I�ҏ m������,�ǏP�� t����3�E�W���� ݟ���:�՟^���[� ��/���S�ܯw� �����8 1߭��� ��w�b�������Z�� ~��ϴ�=�ؿa��� �� �2�D�~������ ��'���K���H߁�� ��@���d��߈ߚ߬� ��G�2�k���*�� N��������1��� U�����N������� n�������Q�� u�4�Xj| �;�_�� ��T�x/� %/���//j/�/ >/�/b/�/�/�/!?�/ E?�/i??�?(?:?L? �?�?�?O�?/O�?SO �?PO�O$O�OHO�OlO �O�O�O�O�OO_:_s_ _�_2_�_V_�_�_�_ o�_9o�_]o�_
oo Vo�o�o�ovo�o�o# �o Y�o}�< �`r���
�C� �g����&�����\��叀�	���-��%�M�ASK 10��'�q��Q�XNO�  `�~���MO�TE  ��!�֑_�CFG ݝ�
��PL_RAN�Gّ?�4���OW_ER 0�R��9�SM_DRYP�RG %0��%�ڏ��X�TART �J���UME_�PROg�y���!�_�EXEC_ENB�  ��5�GScPD͠��$�gTDB2�D�RMS��D�IA_OPTI�ON*�
�7�~��NGVERS������H�I_�AIRPUR(� �ժ��
�F�MT_�Y�TE�ۛ9�OBOT_ISOLC�������K�NAM�E���˿o�_ORD_NUM ?���R��H722  ���������Q�PC_TIMoEOUT*� xQ�oS232��1���C� LTE�ACH PEND�AN������ُ׀Mai�ntenance_ Cons��j���"��ӄNo Usezݶ�|���������"�O�6�NPO��� ����3�C7H_LР	7�#��	��p�!UD�1:��r�RX�VA3IL�����5���_SR  ������~�R_INT7VAL���5�V�����V_DATA_GRP 2���
�� D;�P %���!������� >,bP�t� �����( L:\�p��� ���� //H/6/ l/Z/�/~/�/�/�/�/ �/?�/2? ?V?D?f? h?z?�?�?�?�?�?�? O
O,ORO@OvOdO�O �O�O�O�O�O�O__ <_*_`_N_�_r_�_�_��_�_���$SAF�_DO_PULS�ڐ��o�4�a�PCA)NҚ�4�aF��"�"5}�C�րր
4a���ĵѵ�
Xa�� ���o�o�o �o�o�oyo 2DXVhc�o�r���rXaXad�x�q�q8͑Tesy @�� ����y� ������_ �p.�T���.�k�}�����T D����ŏ׏� ����1�C�U�g�y� ��������ӟ�?�I��y��2�D�	����i�;�oJ��i�pl��
�t��Di��qha~J�� � �g� i�ha`ePaӯ���	� �-�?�Q�c�u����� ����Ͽ����)� ;�M�_�qσϕϧϹ� ��������%�7�I�@[�m�ߑߣߨ��+� ��������&�8�J� \��u������� ������*�/�l�F�0)�������{����� ����������/ ASew���� ���+=O as������ �//'/9/K/��o/ �/�/�/�/�/�/�/�/ ?|�5?G?Y?k?}?�?`�?�?�?0�����p+��0�0�0�0�d`qOO+O=OOO ]GnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o`�o�o�o�o�g��� d'���o,>Pb t������� ��(�:�H�Q�\~�����q�w��M�	12345�678��h!B�!��e���pc � ��$�6� H�Z�l�~������� ˟ݟ���%�7�I� [�m��������ǯح ������1�C�U�g� y���������ӿ���8	��گBH,�T� f�xϊϜϮ������� ����,�>�P�b�t�߫;�j�ߪ߼� ��������(�:�L� ^�p��������D������ �2�D� V�h�z����������� ����
߯@Rd v������� *<N`r1 ������// &/8/J/\/n/�/�/�/ �/�/��/�/?"?4? F?X?j?|?�?�?�?�?@�?�?�?OO&D߆AOSO�/xO�O�O���CB�A��j  W ��h2�b��} �H
�G�/  	ĩB29O _�2_D_V_f\�ogL���1�@3 4 5 6f_�_�_�_�_o o&o8oJo\ono�o�o��o�o�o�o�o�o�^P!r('r-?Qcu �������� �)�;�M�_�q�����B�A g@h@Q�B<��� ��Q  �ɋ㏖�ƂQ>Qt  �@�����`�$SCR�_GRP 1�"X�"al� �� ��� ��E	 j��r���|� hA�������������άM��@�D�` D�@|]��'��ᛊ\R-20�00iC/125�L 567890�PX�PRC2�L g���
V0�5.00 ���� ��vS�H�B��r���@a���a��S�������ǩ	�J�*�<�N��`�h���H��r���v�ѥh�D��y
�-�C3�����ݾĿ�B�r	��������XS����ؾ���@h�ፏh��  @�ȶD����?�XC2#�r�_���%ϠܟIϟ�;ϴEh������BǙ�B�  B�33BƘ��ŗ¨Î�A�@��谘��Ď�@���� ?��ǎ¾@
��ˎ�F@ F�`5� =�4�a�L߅�pߕ߻� �����������.�0�+�=�O�B�]��� ������������!� �E�0�i�T���{_�� �͟������
��t��@+�&��,���R���h1234f�x�F7O��A����� ����Y�� �Q��A �'5J Vh7 ������
/"A�ECL�VL  !���Ѣ�"!L_DE�FAULT*$}��_�uP>#?HOTSTRJ-��"!MIPOWE�RF) �EV%%W7FDOK& V%!"�RVENT 1�1!1!w# L!DUM_EIP/��(�j!AF_�INEJ ?4!�FT�/>>?b?!�a�z?�;�Q?�?!�RPC_MAI�N�?�8��?�?�3V�IS�?�9��?FO!7TP9@PU=O�)�d5O�O!
PMON_PROXY�O��&e�O�OYB�O�-f��O*_!RDM_'SRV+_�)g_v_G!R��_�(he_��_!
�0M�O�,i��_o!RLSY1Nw�*o5g8�_Zo�!ROS�/�l�y4Io�o!
CE[@�MTCOM�o�&k�o�o!	�bCON�S�o�'l�o>!>�bWASRCE_�&�m-�!�bUS	B��(ny�u?� 9S��#�H��l�3��W���'RVICE_KL ?%�+� (%SVC�PRG1����2����3+�0��4�S�X��5{����6�����7˟П򀃤$��9� �_ H����p������ E����m��򁕟� 򁽟8���`��� ���5����^�ؿ� �� ����(��֯P� ���x��&����N� ���v�������� ƿ@�B����҂�ُ 뀋����������� �@�+�d�O���� ����������*�� <�`�K���o������� ������&J5 nY�}���� ��4XjU �y�������/0//T/Ɗ_DE�V �*�M�C:_/q!GRP �2�%� �bx� 	� 
 ,�� 1@K� p� �� � 	� � 2\$�"�" =�$�!� �$�%\#�#����!�!1�!�!\+�#J�� �$1577#p\$�!Y99?  &8-5;C7
8]9�?�# �!%=�?�3�5�!1EO  Q� sa�1�!�%XI�!�$?0w� )�� �!+� 2>OGUt� ]� &� "� *� D�(�$�A�PF!eI�5A9� �$ �9AO�#�!�5�?+[15%5t_�#�(O?;�! 1�!q_?;	5=E�?C7��_"o1�$s� ��0�� �@�    %h-3�#�q��H�8�?
�#� �D1mK?;Ua�8=OkQ1�!�_ S_1	O�oZA~�ew��W���$
�1�v4�o-�� =�c�J���n������� �ȏ����;�"�_��F�X����}	�0X� ��D!uu�  �B� �Rd�a��C7�d �a1A �C7�a�!�o+� �a�a�?W�}�����ʯ ��� ��$��H�/�"�u
T)�3�<�$Yk ���U1�o��u�5�sG�5¯�.8%�?� �!ə-5���W-ϗ�-9 ]����!տ_�A�>�9� b�I߆ߘ�߼ߣ��� �������:�L�3�p� W��{����!��� � ��$��H�/�A�~�e� ��������������  2V=z��� g���
�.@ 'dK�o������//�</I)d� �P�\6��� ���%��2!�A�� ��}M�9U���'lI*g @x��A��3Ai�W�?R�ZA���@1���-������=u����=����%����o�-�?,@����8 @I	r�?�3�@-vy�I)%PALLE�T_HEIGHT�_CHEC�A? �P�	�b%�����z������+�W�B�ӝ¯������V5f!A������o�A��v�@� @<���B��V=­�|��� �.��7Ң²����'V=�N��M>��9�@0@�{�@��)RBZNV9%PLACE_4�LEFTpb�? �P��b%?;+���q�=@�+�K;mW~�F��V>Un�V=�`��>�HFOB��C>(��������CzV=B�3+A������2S�����*N�(�A�x�����7?���q@x;�?W�߰�:�:R1|�?�B,P�&Wb%��R����~��AJ �������u�z�Y�V=@w��&7��B,�V?��0���8@9��*N�W�������e:><-���_e���Z��V=?���A?�q��y��@/���@\4�?%���:PICK�_INCOMING _POIN�O�W!(P�Ji6� ^Bs�B�+=A�¾=\�	A!�MB���>�������
A��#>��H@A�Aɗ��~>�
������>���?du�´�B�7�5�N^1�P?=b����h��%*���$�� ���v_�W�Oof$P����b%�b�������Eu�<�d��,��B4�ɴV=��;��� - @�c5�� �??�A����~>,��A�
�<5��M�}iA����N^��@�`a~��dpA�K��&p��м��?�;?�D��1�P2f!:��m�u ?��� ;Ϭ���#�|���>���{���:@���=;@A���]zERN�(qA�f,��vʷ��1jĜC"���N��/�`���B���>�-K����IA���zGRIPPER_OPEN ?�ogP���b ���" ���f�@H=/�����ؽPl��>����0�A�&���ք��6Β@ICm�V=�4�������ƾ����w$C#���N���X%����?�o�-?�4�� ��v|�QJACKP�O�4��4P���66#������E�������~�fV>��d��7A�	 ?�4�P?�<BAt���~>�c��Q���\[W!¥�
:B�8�>���^R��)��X�ښm@�?'�B<տ�;�? D�)+663��~Bx��B�ͼ�d�A����B�ɉV=>����J�AJ��*��P��+������RN��-�©X��)ͱ� °/\B���>�Ԍ@pٿb>�m�??a:,��iq��^��yg�-7b%B*�\A��s@oP��_�{A��A��q�A�V�AI.A�%��Aڼ@�G����bV>������@���>#�+��Qߍ�B�ʦ>�G����K����f�rg��&2��!��O�L���͔C�b%=?�����t�>��}�<��k�8�O�<e�q�>p����G�A�Um߿Oja�;@�S��XROE�A�������2P^_"��V=�3`�A+_�����@J�@�!��?�����	FI�ND_TOTE �OS,�T�;�<P��Z�b%��i�����@�S�9�:T�%�Vｈ��N��Q���v�A���FA@5�@X4�Pƾ���6���zB�6��0�����A�n�q���0����>?��.@��'�0�KB��T�f� �P�e<�b%���m�l����\ox:�W�~���A�G�٦>���j�JA�h�.�v�J����ƾ���+?K�l����C7Z���������.V>�e]dA^�A��'E�" (@�2�A
������(��e�Zu=��i�-���-e-����=�P���z�{���D��a���b�:A9�@�#�n��+�L��]����ڍ��h +=�*�B�jz�@�1�V����������:;����ks���W���ؔ���hP=����<|B�f2Ij�"���A��q{A����۸IA2����^B�v����>?�_�;�h��¶����Mh�Np��������_��@&'���0a��ϴO��Бv�b ��f!��X�A��$��ɝ�ꒈ���>R�N�����h{B�v?h0�7?�����*N�;�\� rb�<�W�G���c��WC�V>FC��A��������@�Կ ���򙛃\����5P���b%A��a��H���.��f>��-�˟%x���z�"r��@��CA�����h@���A���~>��y����@%��`�2�,�������Nm��bp{��%1A� @�?"�AL�ߚ��;�_̕�4b%:����@B��?�����@?k�;� BQN��h����A����>o0��'<�� ƾ�$@�B�������:�Y|>��!q�@���A��O���%�6s�	�3߿P��eb%<���_?����6�2�?��<圿�;@����AEN�?��?���F��s~>��&@�/���O������¤�B[[�A��`]�@V���^e?�8���!d�NMAI�N IC�5��3�P�jR��e����z=ࡑ��g���o�����N=ք�����A��f?k;�)B�@D�Ŋb�����B���� ~������,�BUKE��,@�>�7��P���@�$F�����;~��D��*�Zu�������@S��@M���z����N{j��m����%��]M�^!��#0f.4�P�A�q?������r��+�A�jT�{B��E��B�������@v�A`h�?0~3�ӱ+��\s?' �����@��n@6��F����@���!�n!���׀	����;�Al�k'�<�M��1��|A��������v�����AJ��A��� ��4�B���BQ@��	?oQBz�^O�>�]�BA�&�a���Am�{��!��=��Ad�h�=�^��~���?*�A�
����@Q�����E޿����Ț���>6�^�j;I���R��nC|��=Ş����X��L���3�>�#:LV_p �fX�RžV]���߀>��I����������~����i/A��Z}�Q�.�@�$Y�f.�@�Akl ����r�LB�@���s0A��V���?V�@�$��I�2_D_*o�1u��֖�ݚBI�N�B�9?�l�>����Ҭ��j=�!���AG���,B�����@k�C�	��s�����.?�����z��`�j��A'A����f����<��y���҄PATH��� �O  P���2R�lU�?�{����:�<�@v ۾	��r��2i���@�����$l@?:R�@.�1Z����M@)����A��@:����SB��O��x�q@Q����ֿ��ņ�R2s�DÅ�/� �խ?��P���Bf ~�A������4��A��B�>�W��r����Aݖ�e@6Β��X����������]�u{���-_����C��j�(��>$���=�s�=���z<�n0���������Aa��)Pz>��)G���Ļ�Y�3>�5^;�+NrΎ`�����A��A>�[p���p����������ܼ>Aì�U����c}�^O����	�@��UU>Z�m�?#�@fk�o��|��O�4P��R���S�rX ?u�4�f�DB�<0�[=���T����&A����?@;3�?7?���H�s���h���~ˡ���K@�^r�����̌Z@��@��������
�H�ֲ)���%��*�%�?\1�;п���Ž���r�*�����5A�`�/?��a@g�%2:?���9�ߩ��~�V2���BBUuj����������@V3�h��݊�oT sK �r�]��F��G���J@��O? (�����?Wo�Z��	����z��[ ���A��ϫ�л�b����Ĉ�d�ֿ)��iy߂BV{���%���)BR3��BU���)`A*wҿpK��0��^%МD��E���j�A �>|�,����i����&�����'>o"�S �@1��?�rS����!�*�6���cD�X�����BY�	Z��DK��_�"B���%�AO�d��A��ظϝ�4�t���]������A���=������¥�)�zN�����������A.�c?���:�^*V�������ɾ��¤�B�����f���ڞ��+�����@$	A��=Y�m�/��(P����u@Գ��3�9��� <�J�����b���7~�c ����6A�>^�9��?��L@i��,f.�9��.��^���������±��B|����P�A����:nA�j7�@�&p?�l��G��$P��ݚF���/��ٻ?,X�������1��O?��JZ�<���3���������lk�����O�8B�����y@�EV|��������^�����kB�NB�"�.B+�~B���
� /.�����5�� �������"[7>8���is�����b>���,�:�30�c�xA�d�?k�f.w��A��n�_���p�S�@�������G��B�l�A�>�����@��Xzߌ�� �. ��5����������S�<�z��L�r������B"���&v��Q,^ґA+a��@`�z� ⿶��aw|�눃� ��^-����B�����.t��=�?%��
GR�IPP����P��
|�u;�f�@(�>����s	?h���;k$�^������?$AL�'���0�WSQ��yږb�W�A5m��~�&�ʡ��q��+U�R~ΐd�n��~�?�����+{��[����/� �P�/�5>��4p����B�S@?���V�?"��Z��Ì������v�A�z!A���@�m1V��z�+�� <��[��g��¿����e9>@�����3�A�����4L��N�����r*�rDk�k=P����5�@`���`B�?��0�3{�����6~?`AA��e?֑A�NA�_�@S�XV��~p��a�����|�������F�`�+Z���|��� �B��������mv�Yy�F?�X?=O|1:�va�q@*l��;s�x;��B	�>��E�Z������h�A�2?/R�Z��P>w������+�=�S���="¦���������J���C�c��������$'f���:V� `TOP:`�/�"I�u=����?���d�S::T@'�߻=�D�ڞ	������A���?!���I�ӿHboV΢�$�@>������8�a�ǤBL�(<~�ę1�����/8��yL�D/��/�_�S��Q���a<�dc�E`�A�ȣ<���[߱w���^<���>@��@
������Af��@Sp6}�4���%?����ɾ�u&|�NC�"s~���W����_²C.t?��9�>���sJACKPO�d�_�b�%P��&��5�yBtEA�����qA���3A��mv����J��A�6�Z�1��_t߁�)/.Z�v]���� �g����?�­>ߚC������A$+&������\��
!�'���Yr*	M�ID_POINT� Pp�:O�rP������w�O����`���A�;�R*���A��ݖ<"�A���@b�:���ґ��3�tB7�q�J3@�V��)"�
���o�A`a�~�0����?$���H��|�_c�P��ö���'�A]E��8�����gA]�OB,c�v��(�ukA��oq?C`����^��Vξ�����'��h7�Q������'�^����@��-
�H����V��2*��j���_�W�P���VE�a���<��!?9�yz��?󲽂C�Z��p�� A�[Ӿ(���@��p@���r_����*�je��T�ߝBL=Fڞ��������O��l>��J0�?���r/�+�o���KVE��z�?���R�tQ�;�O�?R!@����Z�����8�A���h?k�)�ߙ]M��p_B6�)�Aуq����@�Jq�_���ӻ޺��@�>?~������?�AQ�������#��2=����I�u?����:mW~�V��׼��q~������6@t�T�-#�AD��v?����۔��@�����������@�C*|�w~�^8����B�A5d�����@q��>��.���6���!t�|�.�?�[�����������>���?}�A���A���V@�^ٞN$���BVפ��"�Ж��M� ��v�m	�v8�GB�dA��'�f��ܡ��������VE?���?��A�Tx<�A��b+h?at�>�5 �-$A� �l������@��v /B&��BI���v����-�!��"^�%%Ax@0�0U��J+@Z4^��߰��V߁��,P�H�U�N��@��j��7���A�cA=��q^@)����KjA��<�?�\	?���%:��4�!��)�p������qd��P�j`�^?�%%����@א?��PT?2���x!�o�k|S�/�9P�#��]��9T�?�^J��E��ś;�hx~>��K_���Z�����@�����U�U�	������v��Z,���>A��U�L��c����dxB�������%B �A^���CLAMP_CLOSE G �Q�,��P�$�'�	��()^?1�YO��Ƣ�¿����>���b�d�7�;�3�@kq@�>�o"��>�����J�R��O��V�\C�����}����#�B�����/�B"�@������Z����P�A�*V7�bA!7���=�h
�A=�������2��B#$Z=/`��<��_������.�����(7>2���r?����L�����A&���i	����R;��\�ﾫ;P�B�VE��@kAO��@���)>t$ @?�@�ª�E:�2��>pN�A�ec�?���KA����>������U��$.	�r_���+B�s��vQ_+@�Q����N�A��*HB
Yz�$�}�H�D�F�:����@@�������������=��Sm���@? ��@A�0ߖ�Oja���=��@��s��g�Q�fC���>`��~���B�B�f��~�KA���b�tȣ��K"�V@�b���@����[�c��@A�e<����������A��0�������dy�`�>ꎽ�=p�$o���>�>4o��n�����O�>��{�A�AJ\!�������!���3��\���	Ot�Ɵ��k�	��?��)����Y?��H�X4P��%�A�7���@/Ơ�Z�J����BU�1������[Z��h�BN�vN��/��G�?��k��]@*@���@F�;����?�2ߘP�e�VE�1�W��c������y��:���HC?RW5�J� �B���pA�������?3J����C!����1���¾���{¤O���O�5A9}�@�c���`(нSv@>-���K�K�HOME �?�Ou�P�i��be����#T?*J�=��:�R�`���J�b�,p�����A���<��?�0��7���� ���b���E~Z����B�w���@�@75�����3A2�N�@�.]Bl���?���_j�r�j%=��p�A������y;
s	@�i=Y�5B}����� �B���+�{�����/b�*��k��7�>3�M$�q.����M���&A9�D��������uX��%����f���סy�s}���������@�1��5�����t�
G���������6�%�A�ؠA��A��j���������i�?)���g�K���`̮>��{B��8B��� �M��?%_�6�H�~I �P�x��f��p2��0�@�ө)�G^�?�{w�i	�"��Q���V���:R�A�^���v�A��B���3�#*Y���?'��� ���#���{���7�B�����TA�I����&�8|DYt�F�J��@���@!�>�<�?���HB�a�B��o��+�Aۀ�	@AZ}�J$�l������ �����61�?��T�5��C����)b��@�S��&_�'�����&_pA��Y�O ��� @�J�c�����?V=v@p��<���k��1� BY����v@.�@������ۦ@�!Ϝ����z�My�B:,�@)~.���!Í���>���s�B��A��;���kA�#�./��şı��"�����A�ۛ��*����=A���&>�)�{���N
�B8. ?����N��?*�Һ��� �D���e4�xܛ������+�fPA�����G�@�~�Ɓ�+�c
��N|���5P������K���9����p�����p{�=�v����,^���A�-@VrS�>(��v���6��BI�2���@��i�C��l�f������G������ڿV���. @�>#�8m�� �P��A��A�m�V��A�� ��A�n����@�=���������xA�?(@�:�@r�A���xy����m��(�ػ��K���B�gh�^>��yK��?��P����?�1��2�
~Z��THE�_CH�ECKo��P���z��>6��A�Z�?����!���>�?��b����NϲA��G�?�X��&����"��v�3��p�o�K�q@7�����h2]>���A��v�P���V���"����'�~_�<i����P����F���A��?AI�����@�Az�B�<�f������5A�ݞ�?�ք�
���@�1�wʒ��ѝ?䞰���=�·�Q�����^>�~��>�s�F:��?�=���'f�������?�� �P����F�%��A�PAG�ʽ��g@�߅B�Kf�����d�A���@9�����%���YN�!��B��aY��q�ǽ��±W�`BȀ^>��@p�b�8� >y���)���*ck��	M?ID_POI����|h��P��)>5�<�t�����A��(��V��C	�����1���*��A�����@������R���+�*W(���6�1��[���-Ү�����^R���A��@)��@?N1}A.M�V�|����P�"�>5�B���A����A(�}<J���A�z��$���n��J�*�A�O�@��0&����.Bs�Ɓ�
]�?���a<�[·�q!��b�ZN��v>���w�ɡ�O��#@���n������үQe3��19���m?e[J�������@m���=1�o�����[�A�I�@����q����_�R��>2��NK��ISܾ�We�f��iQj�j2<��@�ˡ���g��7��@V3h@���JOGGja��<Q�e:~�����?h��?v���E��>K/u�<�c��.[�I���[1A�����3���P�&�R�����=����3���'�©�x��R@ZN��Ԍ@�q��k������@$�'f@��JR_�SETUPPRO�GRAM��$��Nk~;ň��� �>\�:� ���t���N^>0�c�9A�����Cz@ߓ6Z@�̿�&�H�@��G������`�?�(��-���?�4���c��?��0�J0���������/�N�&&� �з�=�b:"���Ӻ�(��-#���c0�A}����U�U@��S�@��>�&E�@�Љ���+������(�	��W�?���l���X?���d�n9,��C���/�/�?�"�~��a���a�Q�-n�=����:+D/=��`q�x�AŇ5��������D@E��uB?E�@������9���=��(��;���B`@y�T�ZJ@7x�w?�,4����E�?�9G 3"��N�~��]@��s6A D*�������Y��"�DN�WSQ����A�`@�p@��@�&�(���%�g��������u��"�&��:A��><�b?���&�j86��n0fO�?]_��Qf	6
��d�c�T�6?D���#,'�Xߏ��,�N����8�����8X�OA#�����b>��!+������1r>�@ş�U�����-�z�2ө����B�o��� �B�_@~7]CLAMP�� ��3fQf���FJ��������[��< ��+���Ү�����YNA���V!@��{@�6Βz�U�)��h[�������R�£�%��u�ޢL_���ɼ��^k<@���ǿ ���y�(�,oH�f�[~u���=l�ṟ�=��Ү������rA����?�T@"�ϻ?2���^�X����J��>@���U��6��G^�>�,�@A(�u��^����(���8_J[<� �|Qg��$��A׵�A8l����؎A^߫ADL������M{A����=������r��J�ξl5�|��\?�$�B��^¶i_�9�N��OA��+�����?��.t@`5Ͼ����v���>ϯ�!��p�
�
�m���>Nߨ=ט �<-�=�i�=�h0�����A����?�Z}�]zE��c�tl��ӆ?��ѽ�uA�¶���:���>OA����~�@}�d�=��>x�/Њ���}����Z����Va@�˧BX�6��� �����&�yξ��
���?��<B�+0A�p��?�)&�3O���9�}������`�>¤�#���rN��=��h�pA.��@�1��:�ǿ:hu�o�T�  �%�pȲ�jF�����.AsT�<�O���W�3��N{
�o��f���Af��A��A�@AZ�}�4(��6��p�[��g1���Z�����^��E������`0U�#����(�6^?� �TESP�g��ZŽ�QJ��dHG@�0�:�W~��bP�Ϳ5�@�u5����A�\�G�!��@�f�@p����,4�6P��e�e�g�K��~�����G���3L?�'E�w�e�r?:"�B,��D��K�e��Z�=%�����J@� ��;τ�8�y����,B����]MA�*�{���@Iӊ��)��.?P���⎾n�_���^��p������s^>����x?�����e����XA�)"�A�%=��M�<[�4���bM
�v��ZA�,:����<A���µ�y�{��@0L�.ߘ¹�Q�9�����?v@�7���P����@d6ſ�]�����+��������^H`�w��=&���i!�@(��^!�~}@��A��िOja@�� A�P�Pr����>+�����^�´Z���1g�������W��+��@�ņ�F/�����w��HO�ME ��z�u�����T�����z��Ԍ_>9lZ�����;Z��^�a��D5��A��H��7�ަQ@��^�/�3��}��]���d�A¬��}�����$c�*��&��-s��@N�q��;_��%�V� !eG_CH�qK���������*����+�=�J��~������^�[�	�E�5A��5���ݰ@���@��x�^����������������+��7
���D'�/ �J\�!@R���z<�����b�ER�_OPEND�V�$��A�4;�����,�=XS����s�Q1���^G�@��A��L��h�@��y@���j�b�8/���^���옾�\;¦������
���-$���e�i���@;_̊2Is�
 q�X�=����6}A��iA�Ks���A-�>���F.��P���zA����@�+��C���@���B4����#g�;�׾r²�ߛ���
�i@��A#�g����H��7�@�+��s����������Y:���@?�zA�7=������?����
���L�ڻ+�A��b����@���M�e�
�C+�&�2����m ��M���³/���m.�I|@�J�3Y�?�� v;?�����HT  #P���jž�I�@�� �E�����V�Bb��>�!�
�����B,�'@S���[���^�.���./�.�ھi�L��<����_$P�J[�nY@��0��"����9*�MAI P?LASTICi���  P�8<��~A����b�<_`A��m�=�.�ޮ�����`@BJ�;��$��ڼ�/�@�����;�&���C�>0R�¿x(���I����yKA��7���S���4_����
����INCOM�br?GE_;P�I���2��t@����d��V�@U��<���Op�$ؿFA���?��r/>��vޮ�����ø���l^>@���W^q��b
�����A����=aj�٠���(\�8V"O�4G&a_R5B`a��$SERV_\0LW  :uHP�Aa>2TOUTPUA@?V_B`@2T�RV 2���q� � ("si�p�>�pb  3�q]�2TSAV&``ZLYTOP10 2~Y� d � \�� p  �J`2C`e� sB`Ƃ�P�U�B`>J`B`�iP�qJ`�2c�d�*`
�Vohozo�o �o�o�o�o�o�o
 .@Rdv��� ������*�<� N�`�r���������̏0ޏ����UYP�_NS�FZN_CFG y&KSTmQ|�U8�GRP 2�F��Q ,B �  A���QD;�� B���  B�4SRB21ޱVHELL;� 
��V�P�P\Y����RSR����� F�1�j�U���y����� ���ӯ���0��T��e��Q�\�  �:a%e�����s�s���Q*`�����޽���	`�Pm�����HK 1�� (bÿ`Ϧ^{ύ϶ϱ� ����������F�A߀S�eߎ߉ߛ߭ߩ�OMM ���߬��FTOV_ENB�=T:a�U;�OW_R�EG_UI�ORIMIOFWDL����ޅ�P�WAIT���Z�x�XP<�܅Tu�TIM<������VA<P��P�_�UNIT����YL]C5�TRY<��U��PMB_HDD�N 2~[  (`��a�W� x��s� ���������������$8�ON_ALI�AS ?)&iS( he�QZl~�� �V����) ;M_q��� ���//%/7/I/ �m//�/�/N/�/�/ �/�/?�/3?E?W?i? {?&?�?�?�?�?�?�? OO/OAOSO�?wO�O �O�OXO�O�O�O__ �O=_O_a_s_�_0_�_ �_�_�_�_�_o'o9o Ko�_\o�o�o�o�obo �o�o�o#�oGY k}�:���� ���1�C�U� �y� ��������l����	� �-�؏Q�c�u����� D���ϟ�󟞟�)� ;�M�_�
��������� ˯v����%�7�� [�m������N�ǿٿ �����!�3�E�W�i� ύϟϱ����π��� ��/�A���e�w߉� ��F߬��������� +�=�O�a�s���� ���������'�9� K���o�������P��� ��������5GY�k}��$SMO�N_DEFPRO�G &����� &�*SYSTEM*���@+ �R�ECALL ?}��	 ( �}3�xcopy fr�:\*.* vi�rt:\tmpb�ack=>10�.$202.21:19680 2�;M_o}4a�/8��� �}8s:ord�erfil.da�t���J/\/n/}=/mdb:�'/ 43/�/�/�/{� &�/I?[?m?�?#? ��?�?�?�/�/�/ EOWOiO|/�/)O�/�O �O�O�/�?�?0?A_S_ e_x?�?_�?�_�_�_ �?O�O,O=oOoaotO �O!o�O�o�o�o�O_ �_(_�oK]�o�_ %8��� oo�o �oG�Y�k�~o��o4� ŏ׏��o��2C� U�g�z�����ӟ ��
���.�?�Q�c� v���#�����ϯ�� ���*�;�M�_�r�������:�˿ݿp�x�yzrate 124 ������D�V��h�{��#�8:172�"�4��������� �ϡϳ�D�V�h��{�!��69.25�4.14&�4:16120 %�7���������tpdisc 0�ߠҢߴ�E��W�i�|�tpconn 0�� �2�������z�:��� ��=�O�a�t�1���@��6�������~�5��͡����K]��6��& :��p ������I[m�� �6������ �4E/W/i/|// ��/�/�/��0 A?S?e?x�%?��? �?�?�/�/,/=OOO aOt/�/O�/<O�O�O��L�$SNPX_�ASG 2����Q�7  �B%��O6_�  ?��FPAR�AM U^Q �	$[P9T�� 9X�T��PPOFT_KB_CFG  �#�U�COPIN_S_IM  [�R��_�_ocPRV�NORDY_DO�  �U�U#bQSTP_DSB�^��Rgo�KSR �Y � & �PNS0001� PROGXQEI�GHT_CHEC�K�Ysd�STOP_ON_ERR0o��B�aPTN zUp�A�b�RING_PRM��oBbVCNT_GOP 2 U�QPx 	�V�YePs|}�ZPr��p��t��w�JVD7pRP 1!^Y�Pvqa� ����0�W�T�f� x���������ҏ��� ��,�>�P�b�t��� ������������ (�:�L�^�p������� ��ʯܯ� ��$�6� H�o�l�~�������ƿ ؿ����5�2�D�V� h�zόϞϰ������� ��
��.�@�R�d�v� �ߚ��߾�������� �*�<�N�`���� �����������&� M�J�\�n��������� ������"4F Xj|����� ��0BTf x������� //,/>/e/b/t/�/�/�/�/�rPRG_�COUNT�V�r�)ENB�%M�3�T?_UPD �1"�kT  
 �/|Bd?v?�?�?�?�? �?�?�?OOAO<ONO `O�O�O�O�O�O�O�O �O__&_8_a_\_n_ �_�_�_�_�_�_�_�_ o9o4oFoXo�o|o�o �o�o�o�o�o 0YTfx��� �����1�,�>� P�y�t���������Ώ ��	���(�Q�L�^� p����������ܟ�  �)�$�6�H�q�l�~� ������Ưد������,_INFO 1=#R580Z�	 1�u�`�����<���(���ÿ����཭��������뾻���¤@k�፥�|��� D��z�?��C2��ݗ边��DB�&�8�� Y?SDEBUG� S0��(�d;9c�SP_�PASS�%B?~u�LOG $O�]\1  (����?��(�.�  ��71(�
MC:�\�Ģ��)��_MPC�� ����.���/UD1��25��?SAV %��1����*�Q�SV�b�TEM_TIM�E 1&��]0� 0 ��'���� 4�*�4��Fc4�p���MEM�BK  R571�����7�I�Y�X�|80� @Y�&���{���t���������@���)� ;�M���f�x����������� �����
�.@Rdv��,e �����( :L^p�������� //��SK ���!"�R/d/v/j�;�80  x/���/62&�$����/�)=(���!O�*��C=PC?_65>c�g� �?d?�?�?�?���?�,�O9OKO]OoO�O(�$�O�O��O�O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_�_o#o�/T1SVGUNwSPD�� 'u���F`2MODE_?LIM '��y�2Bd2O`oa(��Ae�ASK_OPTI�ONj��y��a_�DI��ENB  ���u��aBC2_?GRP 2)5%u�0����@C�"s:l�BCCFG +��k(��2*�Yz` w�������	� �-��Q�<�u�`�r� ����Ϗ���ޏ�� '�M�8�q�\������� ��ݟ���ڜ	�۟<� N�ɟ+���o�����̯ ڪ5%�������� >�,�b�P���t����� ���ο��(��L� :�\ς�pϦϔ��ϸ� ������ ��H�.�� \�nߌߞ߰�.����� ��
���.�@�R� �v� d����������� ��<�*�`�N���r� ������������& 68J�n�Z� �����4" DjX����� ���//./0/B/ x/f/�/�/�/�/�/�/ �/??>?,?b?P?�? t?�?�?�?�?�?O� O.OLO^OpO�?�O�O �O�O�O�O __�O6_ $_Z_H_~_l_�_�_�_ �_�_�_�_ ooDo2o Tozoho�o�o�o�o�o �o�o�o
@.dO |����N�� �*��N�`�r�@��� ������ޏ̏���� 8�&�\�J���n����� ��ڟȟ���"��F� 4�V�X�j�����įz ܯ���0���T�B� d���x�����ҿ���� ���>�,�N�P�b� �φϼϪ�������� �:�(�^�L߂�pߦ� �߶߸��� ���$�گ <�N�l�~����� ������� �2� �V� D�z�h����������� ����
@.dR t������ �*`N�:� �����n//�$/J/8/n/X&� �$�TBCSG_GR�P 2,X%��  �� � 
 ?�   �/�/�/�/�*�� ? ">?E?/?i?{=�"�#�.�,d����1?�!	 HC�; {6&ff�2� �{5�1A��!�?�9Dw)�{6��F�|4AB4�?�?HL�@YA�8$B�:O�MCwj��PN333{5?B�C�O�O��O{9�O_�N|4>�LG�AB�_Z]@�8 [6�8�U�_^_p_�_�_@�_�_o#o2kh�La	V3.002b�	rc2l2c	�*n`fd�"}o<fG��?�33� X��ai �`�m�o � �# _�o�e�!J�2�#/�-�o
xC�FG 1X%X�!�!4z��"�b94�x��� �za �����+� �O�:�s�^�p����� ͏���܏� �%�K� 6�o�Z���~�����۟ Ɵ؟���5� �Y�k� q��v�����D�ͯ�� ݯ��'��K�6�o� ������`�ɿ���ؿ ��#ό!x/H�T/X�Z� lϢϐ��ϴ������ ���D�2�h�Vߌ�z� �ߞ�������
���.� �R�@�v�d���� ��������0��� P�r�`����������� ����&8��HJ \������� �4"DFX� |������
/ 0//T/B/x/f/�/�/ �/�/�/�/�/??>? ,?b?P?r?�?B��?�? �?~?O�?OO(O^O LO�OpO�O�O�O�O�O  _�O$__4_Z_l_~_ 8_�_�_�_�_�_�_�_  oo0o2oDozoho�o �o�o�o�o�o�o
 @.dR�v�� �����*�<��? T�f�$�"�����̏�� ��ޏ ���J�\�n� ,�~�����ȟ����� �"�ܟF�4�j�X�z� ����į���֯��� ��0�f�T���x��� ��ҿ������,�� P�>�t�bτφϘ��� H�����
ߴ�:�(�J� p�^ߔ߂߸ߦ�����  ����6�$�Z�H�j� ����n������� ��2� �V�D�f���z� ������������
 R@vd��� ����<* `rߊ�"�X� �/�&//6/\/J/ �/�/�/b/t/�/�/�/ �/"?4?F?X??|?j? �?�?�?�?�?�?�?O OBO0OROxOfO�O�O �O�O�O�O�O�O_>_ ,_b_P_�_t_�_�_�_ �_�_o~�.o@o�_ o^opo�o�o�o�o�o �o$6HlZ |~������  ��D�2�h�V�x�z� �����ԏ
���.� �>�d�R���v����� П�������*��N� <�r�`�����Ro��ү 䯎���8�&�H�J� \�������ȿڿ쿪�����4�"�X�B�  9~��� �Ɩ�����$TBJOP_GRP 22J���  �?���	�µ�4����R� ��� �,�^�� ��� � s � ���� @~���	� �C� 2�Q?p�D������N�&ffV�K�W�i��<9]2�?�ߚ?L�͊�BH�  A�Hץ߰�D�)���>��SBF�Y����g��� �����>���<�����?333?f�h��B�  B x��=���D5mF���n�w�ы��Af�����C+�&�.���Cj�����߁�����;ć�B����Ⴔ����]���������<w��6����F� ��j�|�N�O��"(�8���z�J6����>���C4(� ��}����� ���&@*\ f�r�����(�'/����ưJ!N�	V3.00���rc2l��*�t ��}��/�' �F�  F�  �GX G7� �GR� Gr0 �G�� G�@ �G�� G�\ �G�� G�` �G�� H
� �Hd H" �H.� H;� HH2 HUޝ"�E�� E� �!F�@ F� Fj`� F�� F�� �"�!� G$w G� GVص#��� G�L G��� G�h G��� =u=�+,XZ5�Ќ�r?�2���3?��  &����ESTPAR v������HR�0ABLE ;15�� �0�0RDD����|:
�'�(�(�ǉ��'	�(
�(�(A��U�(�(�(�6'RDI�?���FA�����7OIO[OmH�DO �O�K�O_ _2_D^�2	S�O�� �Joo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [���P�_��C�}�_ �_�_�_gOyO�O�O�O��H�2�rNUM  �J���"��� @�@�2_CF�G 6k��&�@���IMEBF_T�T�1����0��VE�R�CAÆ��R {17K 8/f�� ��P�
 M��  ���*�*�)� ;�M�_�q��������� ˟ݟ���\�7�I� ��m��������ǯٯ|���  PDT�&� � "[L�^� �C{�M!�����UK�8��ѿ�_DE��ώ �OTF,�>� �c$Cd�v� �$��ϲ���s�����R#ID���_e�چ�@��0MI_CWHAN�� � �ӿDBGLVL�����1��ETHER_AD ?�5��m��00��:e���4:71:d0:�66 ��7��68��69��ROUT6׀!iZ!<�Z���9��SNMASK������255�.��2.`#���5������0OOLOF/S_DI Tռ��ORQCTRL C8��PS�?8�T'� \�n������������� ����"4FXj�|�K�����2P�E)�TAI����P�GL_CONFI�G >k�{����/cell/$�CID$/grp1�M_q��KS������// �>/P/b/t/�/�/'/ �/�/�/�/??�/�/ L?^?p?�?�?�?5?�? �?�? OO$O�?HOZO lO~O�O�O1OCO�O�O �O_ _2_�~}�Oh_ z_�_�_�_�_0���_�]��Oo1oCoUogo yo�O�o�o�o�o�o�o �o-?Qcu� ������� )�;�M�_�q������ ��ˏݏ�����7� I�[�m���� ���ǟ ٟ������3�E�W� i�{�����.�ïկ� ������A�S�e�w� ����*���ѿ������+�&�Us�er View �;}}1234567890\�nππ�Ϥ϶Ͼ�G�����B�2Oɻ� �2�D�@V�h�z�����I�3� ���������"��C���4��|��������5�����5k�0�B��T�f�x��������6 �����,>��_��7������ ��Q��8�L ^p������ lCameraM�C// 0/B/T/f/DRE��/ �/�.Z��/�/�/??(?�  ���x? �?�?�?�?�?y/�?O Oe?>OPObOtO�O�O�����/O�O�O_ _,_>_�?b_t_�_�O �_�_�_�_�_o�O�G j�_Poboto�o�o�o Q_�o�o�o=o(: L^po�GD;	� ������o<�N� `����������̏ޏ ����s�(�:�L�^� p���)�����ʟ��  ��$�6�H�G�	 ߟ������ʯܯ� �$�6���Z�l�~��� ����[��G:K� �� $�6�H�Z��~ϐϢ� ���������� �ǿٷ9��a�s߅ߗߩ� ��b��������9�@K�]�o���"	�0���������(� ��L�^�p������� ������������� GYk}��H�� ��41CU g�[;���� ��/�1/C/U/� y/�/�/�/�/�/z�� �Kj/?1?C?U?g?y?  /�?�?�??�?�?	O O-O?O�/�%3k�?�O �O�O�O�O�O�?	__ -_xOQ_c_u_�_�_�_ RO�%�{B_�_	oo-o ?oQo�Ouo�o�o�_�o �o�o�o�_�%� �ocu����do ���P)�;�M�_�xq���*}  .y ��ď֏�����0��B�T�f�x�   �C��o�2o�D���?�-�B�  C3��*q��ɺ�����*q@+� BS���h�[*p?�łBl@֑v������z�ǟ Aǒ�^"�\��x6FB o�Ο\�������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ���ϲ�������&� 
�*p(  覀( 	 ��0��T� B�x�fߜߊ߬߮���@������>�,��� ������� ��������%�,sr� O�a�s���������� ����8�'9��] o�������� �F#5GYk} ������/ /1/C/U/�y/�/�/ ��/�/�/�/	??b/ ??Q?c?�/�?�?�?�? �?�?(?:?O)O;O�? _OqO�O�O�O�O O�O �O_HO%_7_I_[_m_ _�O�_�_�__�_�_ o!o3oEo�_�_{o�o �o�_�o�o�o�o doASe�o��� ���*��+�r O�a�s��������� ߏ��J�'�9�K�]� o���ȏ����ɟ�� ���#�5�G���k�}� ��֟��ůׯ����T�4�@ /�<�N��`�/�6����)�frh:\tpg�l\robots�\r2000ic���_125l.xml�Ŀֿ������0�B�T�f�r��� rϗϩϻ�������� �'�9�K�]�t�nߓ� �߷����������#� 5�G�Y�p�j���� ����������1�C� U�l�f����������� ����	-?Qh� b������� );Md^� ������// %/7/I/`Z//�/�/ �/�/�/�/�/?!?3?�E?W>y��� |6���<< �� ?�W;�?W?�?�? �?�?�?O�?0ONO4O FOhO�O|O�O�O�O�O�_�O�O_J_X���$TPGL_OUTPUT Ab��b� z0��x6FB�PZR�?łB4  �Qb����ɺ�����ZR5/�B�  �1��^��_�_�_ oo)o;oMo_oqo�o �o�o�o�o�o�o�%7Ewz0�OPce�ll/cont1�/grp1/dc�s/cpcz/z�6/f �eB��� �,kB�P�X��q ���gB^����X�7��@^���� �QBО�X�t�u^��p�XO�rH�u[mx1y�u��p��q�ZOBX��s$A�r�u��֊s�<���v2345678901f�x��� ������ȃ�sd���� �&�8�J��s}M�u� ��������U�g��� �)�;�M��[����� ����˯c�ٯ��%� 7�I���������� ǿٿq���!�3�E� W��eύϟϱ����� m����/�A�S�e� ��sߛ߭߿�����{� ���+�=�O�a���� �������������@'�9�K�]�o�׍}u1�������������
@�|?.@�: ( 	 Cuc�� ������; )_M�q��� ��/�%//I/7/�Y/[/m/�/�/�/Qv� x0�6�/?=�/5?G? !?k?}?Kz�/�?�?Z? �?�?�?�?,O>O�?BO tOO`O�O�O�O�O�O PO�O(_�O_^_p_J_ �_�__�_�_�_�_o $o�_0oZo�_�_�o�o <o�o�o�o�o ~o DV�oB�fx� �2�
���@�R� ,�v����p���Џj� �����<���$�r� ������������N� `�&�8�ҟD�n�H�Z� �������쯆�د"� 4��X�j�ȯR���:� ��ֿ�¿��|�� T�f� ϊϜ�vϨ��� 0�B��ߴ�"�P�*� <߆ߘ��ϼ���hߺ�������:�L��")�WGL1.XML�
���$TPOF?F_LIM � ��!���Nw_SV��  ���P_MON �B�%�����2��STRTC�HK C�%�������VTCOMP�AT��H��VWV_AR D��k�.�� � �� �����_DEFPROG %��%  R_SE7TUP��RA�������_DISPLA�Y�����INST�_MSK  � ��INUSE9R>���LCKG�QUICKMEN�k��SCRE� ��%I�tps�c��G� �	�� _�	ST<���RAC�E_CFG E���k���	��
�?�HNL 2!F��� *r� ��^ p��������ITEM 2G�J �%$12�34567890<1/C%  =<;/a/<s/{#  !�/�+��E/�/��//�/S/ ?%?�/;?�/�/�?�/ �??�?�?_?O?a?s? �?�?O�?gO�O�OO �O'O9OKO�OoO_A_ S_�O__�O�O�O�_�_ 5_�_ok_o�_�_jo �_�o�_�o�oo�oCo �oyo9�oIo� �o�	-�Q� #�5��Y����e� }��׏�M���q��� L���g�ˏ������� %�7� �[���+�Q� ןǟٟ�����3� ߯��{�;�����ï =�篓���˿/�׿S� e�w���Iϭ�m��� ������=���a�!� 3ߗ�I߻�ߖ��ϱ� �������]��ߓ� �����u������ 5�G�Y������O�a� ��m����������C� y�+����x�SH}
� 3 �}
 "���
 ��+~�
UD1:\8����R_GRP� 1I+� 	 @��@�������  $/2*�8\/G/�/k%?�  �/�+�/�/ �/�/�/??%?'?9? o?]?�?�?�?�?�?�?�?O	K%O7O��SCB 2J� �/�O�O�O�O�O��O�O__�UTORIAL K��^_�V_CON?FIG L��z��_n\OUT?PUT M�	�P���_oo1o CoUogoyo�o�o�o�o��o�o�Q�\Re�gular Option�o0B Tfx����������_�!�3�E� W�i�{�������ÏՏ ��d��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� �������������U����_9K]o� ������� �5GYk}�� �����/1/ C/U/g/y/�/�/�/�/ �/�/�/	??,/??Q? c?u?�?�?�?�?�?�? �?OO(?;OMO_OqO �O�O�O�O�O�O�O_ _$O7_I_[_m__�_ �_�_�_�_�_�_o!o 2_EoWoio{o�o�o�o �o�o�o�o.oA Sew����� ����*=�O�a� s���������͏ߏ� ��'�8�K�]�o��� ������ɟ۟����#��C�B�J��X�>�-��"\R�egular Option����ί ����(�:�L�^� p���5�������ѿ� ����+�=�O�a�s� ��6��ϻ�������� �'�9�K�]�o߁ߒ� �߷����������#� 5�G�Y�k�}��߳� ����������1�C� U�g�y���������� ����	-?Qc u�������� );M_q� ������// %/7/I/[/m//�/� �/�/�/�/�/?!?3? E?W?i?{?�?�/�?�? �?�?�?OO/OAOSO�eOwO�O�O�$TX�_SCREEN �1NV�>��}��O�O�O__(_:_�O���Oz_ �_�_�_�_�_K_]_
o o.o@oRodo�_�o�_ �o�o�o�o�o}o* �oN`r��� 1����&�8�� \����������ȏڏ Q���u�"�4�F�X�j� |�����ğ֟��� ���0���T�f�x���𜯮�%�ү�$UA�LRM_MSG k?�I��@ ʯ �:��G�:�k�^��� ���������ܿ� ��1��SEV  ��c��ECFoG P�E�A�  �5@�  }A��   BȦ2�Q�@�����l� �A �Qg�ª�Gu4P�������nP�3�����ą�A�Yx�Qe<'��TyQ�e�
��_Qf� $"��0Qf�L��Y{Qf��:�X�Qf�!� ��NQf�o�G�RP 2Qy� 90�¦1	 2�����I_BBL_N�OTE Ry�T��l�2��@�1����DEF�PRO�%� �(%CLEAR�_IO LOSE� CHECK T_J�7:�l�W�%Ϝ� ������������,��>�)�b���FKEYDATA 1S�I���p �ǟ6�����������
��,�(=�4(PO?INT  ]EG  OON����tNDIRECT�<�I�OICE`��TOUCHUP���� RE INFk�#`rY�} �����/&//�J/1/n/�/�����/frh/gui�/whiteho?me.png�/�/��/�/�/?��&point�/<?N?`?�r?�?6  �%look+2�3�?�?�?�?� O�?�6indirec*?FOXOjO|O�O�>clos�$9O�O��O�O__0�&t?ouchup6ON_�`_r_�_�_4�&arwrg5O�_�_�_ oo�H5oGoYoko}o �o�o0o�o�o�o�o �oCUgy�� ,����	��-� �Q�c�u�������:� Ϗ����)���M� _�q����������%�� ���	��-�?�F�c� u���������L��� ��)�;�ʯM�q��� ������˿Z���� %�7�I�ؿm�ϑϣ� ����V������!�3� E�W���{ߍߟ߱��� ��d�����/�A�S� ��e��������� r���+�=�O�a��� ������������n��� '9K]o���@������+��� �4F�""o��#,g/�_(OINT  ]��� IRECT <��  ND�/�/ CHOICE��:/�UCHUP e/f/�/�/�/�/�/�/ ?�/3??W?i?P?�?�t?�?�?�?�?Ɲ&Ewhitehom�D� O2ODOVOhOw�Fpoin�_�O�O�O�O��O�Oi/direc�O0_B_T_f_x__/in_�_�_�_�_x�_�_�AclosD��_>oPoboto�o�Jt?ouchup�_�o��o�o�o�Narwrg�_@Rdv� ������� *�<�N�`�r�����%� ��̏ޏ������8� J�\�n�����!���ȟ ڟ����"���F�X� j�|�����/�į֯� �����?��T�f�x� ��������ҿ���� �,ϻ�P�b�tφϘ� �ϼ�K�������(� :���^�p߂ߔߦ߸� G����� ��$�6�H� ��l�~������U� ����� �2�D���h� z�����������c��� 
.@R��v� ����_� *<N`���� ���m//&/8/hJ/\/3�j+�@j/�/�/B�/�/�/� C,�??�8OIN�T  ]%?'? I�RECT Q?R? � NDf2}?? CHOICE@?�?80UCHUP�?�?O %OOIO0OmOOfO�O �O�O�O�O�O�O!_3_�_W_6��Uwhitehom&d�_�_�_��_�_��fpoin�/o-o?oQoco�_i?/direc
o�o�o�o�o�owo/in �o!3EWi�oachoic�_������/touchup�.�@�R��d�v��^arwrg ��ԏ����� .�@�R�d�v������ ��П������*�<� N�`�r��������̯ ޯ����&�8�J�\� n�����!���ȿڿ� ��ϟ�4�F�X�j�|� ��e_+���������� �%�B�T�f�xߊߜ� +�����������,� ��P�b�t����9� ��������(���L� ^�p���������G��� �� $6��Zl ~���C���  2D�hz� ���Q��
// ./@/�d/v/�/�/�/ �/�/_/�/??*?<? N?�/r?�?�?�?�?�?ڣ��;�sP���OO'M�?IO[O5F,G_�O?_�O�O �O�O�O
_�O._@_'_ d_K_�_�_�_�_�_�_ �_�_o�_<o#o`oro Yo�o}o�o�o���o &8JY?n�� ����i��"� 4�F�X��|������� ď֏e�����0�B� T�f�����������ҟ �s���,�>�P�b� 񟆯������ί�� ���(�:�L�^�p��� ������ʿܿ�}�� $�6�H�Z�l�~�Ϣ� ���������ϋ� �2� D�V�h�z�	ߞ߰��� ������
��o.�@�R� d�v��߬������ ������<�N�`�r� ����%��������� ��8J\n�� �3����" �FXj|��/ ����//0/� T/f/x/�/�/�/=/�/ �/�/??,?�/P?b? t?�?�?�?�?K?�?�? OO(O:O�?^OpO�O �O�O�OGO�O�O __�$_6_H_�J[�>����s_�_ �]o_�_�_�V,�o�_ �o ooDoVo=ozoao �o�o�o�o�o�o
�o .RdK�o� ������*�<� �`�r����������O ޏ����&�8�J�ُ n���������ȟW�� ���"�4�F�՟j�|� ������į֯e���� �0�B�T��x����� ����ҿa�����,� >�P�b��ϘϪϼ� ����o���(�:�L� ^��ςߔߦ߸����� ��}��$�6�H�Z�l� �ߐ���������y� � �2�D�V�h�z�Q� �������������� .@Rdv�� �����*< N`r���� ��//�8/J/\/ n/�/�/!/�/�/�/�/ �/?�/4?F?X?j?|? �?�?/?�?�?�?�?O O�?BOTOfOxO�O�O +O�O�O�O�O__,_ �OP_b_t_�_�_�_9_ �_�_�_oo(o�_Lo�^opo�o�o�o�o����k�������o�o}�o);v,'�l��w�� ���� ��D�+� h�z�a�����ԏ�� ��ߏ��@�R�9�v� ]�������П���� �*�9oN�`�r����� ����I�ޯ���&� 8�ǯ\�n��������� E�ڿ����"�4�F� տj�|ώϠϲ���S� ������0�B���f� xߊߜ߮�����a��� ��,�>�P���t�� ������]����� (�:�L�^�������� ������k� $6 HZ��~���� ���� 2DV ho������ ��/./@/R/d/v/ /�/�/�/�/�/�/�/ ?*?<?N?`?r?�?? �?�?�?�?�?O�?&O 8OJO\OnO�OO�O�O �O�O�O�O_�O4_F_ X_j_|_�__�_�_�_ �_�_o�_0oBoTofo xo�o�o+o�o�o�o�o �o>Pbt� �'�������(�� *��� ���S�e�w�O�������,��܏�� � �$�6��Z�A�~��� w�����؟�џ��� 2�D�+�h�O���s��� ¯���ͯ
���@� R�d�v��������п �����*Ϲ�N�`� rτϖϨ�7������� ��&ߵ�J�\�n߀� �ߤ߶�E�������� "�4���X�j�|��� ��A���������0� B���f�x��������� O�����,>�� bt�����] �(:L�p �����Y� / /$/6/H/Z/1�~/�/ �/�/�/�/��/? ? 2?D?V?h?�/�?�?�? �?�?�?u?
OO.O@O ROdO�?�O�O�O�O�O �O�O�O_*_<_N_`_ r__�_�_�_�_�_�_ _o&o8oJo\ono�o o�o�o�o�o�o�o�o "4FXj|� �������0� B�T�f�x�������� ҏ������,�>�P��b�t�����o ��}�o ���ß@՟睿�	����,� L���p�W�������ʯ ��� ��$��H�Z� A�~�e�������ؿ�� ��� �2��V�=�z� ��k/����������
� �.�@�R�d�v߈ߚ� )߾���������� <�N�`�r���%�� ��������&���J� \�n�������3����� ����"��FXj |���A��� 0�Tfx� ��=���// ,/>/�b/t/�/�/�/ �/K/�/�/??(?:? �/^?p?�?�?�?�?�? ���? OO$O6OHOO? lO~O�O�O�O�O�OgO �O_ _2_D_V_�Oz_ �_�_�_�_�_c_�_
o o.o@oRodo�_�o�o �o�o�o�oqo* <N`�o���� ����&�8�J� \�n��������ȏڏ �{��"�4�F�X�j� |������ğ֟��� ���0�B�T�f�x�� ������ү�����0�
���0���3�E�W�/�y���e�,wϼ�o��ǿ� ���:�!�^�p�Wϔ� {ϸ��ϱ������$� �H�/�l�Sߐߢ߉� �߭������? �2�D� V�h�z������� ����
���.�@�R�d� v�������������� ��*<N`r� �%���� �8J\n��! �����/"/� F/X/j/|/�/�///�/ �/�/�/??�/B?T? f?x?�?�?�?=?�?�? �?OO,O�?PObOtO �O�O�O9O�O�O�O_ _(_:_�^_p_�_�_ �_�_�O�_�_ oo$o 6oHo�_lo~o�o�o�o �oUo�o�o 2D �ohz����� c�
��.�@�R�� v���������Џ_�� ��*�<�N�`�� ������̟ޟm��� &�8�J�\�럀����� ��ȯگ�{��"�4� F�X�j���������Ŀ ֿ�w���0�B�T��f�x��$UI_I�NUSER  ������?�  y�}��_MENHIST� 1T��_  (��QP�(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,181,�1 �17 VERIFY�)�;�M��_��'���34,�4 1 ALIB�RATION� EFT'�����d�v���7�TUPPR�OGRAM�ET,22 H��G�Y�������4��LAS�TIC_PALLET_L��8���������Ϗ�148,2�  ��HEIGHT_CHECK7�`Q�c�����53�@��4���������)�����13��ACKPO��00 ��Ug�y|�,70FP����������� ���.@Rdv� ���� �/�+/=/O/a/s/ �//�/�/�/�/�/? ?�/9?K?]?o?�?�? "?�?�?�?�?�?O�? 5OGOYOkO}O�O�O0O �O�O�O�O__
C_ U_g_y_�_�_�_�O�_ �_�_	oo-o�_Qoco uo�o�o�o:o�o�o�o );�o_q� ���H���� %�7��[�m������ ��ǏV�����!�3� E�0_N�{�������ß ՟؏����/�A�S� �w���������ѯ`� ���+�=�O�a�� ��������Ϳ߿n�� �'�9�K�]��nϓ� �Ϸ�������|��#� 5�G�Y�k�V�ߡ߳� �����������1�C� U�g�y�������� ����	���-�?�Q�c� u�������������� ��);M_q� �$���� �7I[m�|���$UI_PAN�EDATA 1V������  	�}c�/frh/cgt�p/flexde�v.stm?_w�idth=0&_�height=1�0��ice=T�P&_lines�=15&_col�umns=4�f�ont=24&_�page=who�le��z�)p�rimA/j/  }�m/�/�/�/�/�/�/ )�/?�/5??Y?k? R?�?v?�?�?�?�?�?�OOOCOz���� c@ ���{$���2�
%3�@.1(%do�ub�@2MO+Hua�l�O
_qKitree�A_E_W_i_{_�O �_�_�_�_�_�_o�_ /ooSoeoLo�opo�o�o�o�oVH � �c@	 "�0�sO�O�OP3
&( ��O(%t#p3�o�khird��~/�� ���)��oM�4�q� ��j�����ˏ��ݏ� �%��I�[�B���o�q 	2W�. t��ǟٟ����b� !�E��i�{������� ï*��ί����A� (�e�w�^�������ѿ@����ܿ�+��bB� �_�d�vψϚϬϾ� ���U���*�<�N� `��τߖ�}ߺߡ��� �������8��\�n� U��y����;�M��� �"�4�F�X���|��� ������������s� 0T;x�q� �����,> %b������� ��E/(/��L/^/ p/�/�/�//�/�/�/  ?�/$??H?Z?A?~? e?�?�?�?�?�?�?o �?/DOVOhOzO�O�O �?�O5/�O�O
__._ @_�Od_v_]_�_�_�_ �_�_�_�_o�_<oNo�5oroYo�o�oO-D���o�o�o
.@) �oe�ET���� ��R��3��,� i�P���t���Ï��� Ώ���A��H+C%K��$UI_POSTYPE  +E�� 	 �`�� �����C�s�QUICKME�N  �� �����_RESTO�RE 1W+E����*default�K�  INGLE~�PRIM��momenup�age,1388,1,27N���������� m  d�290,1����� '�ʦB�T�f�x����� 4�����/��
� �.�@�R���vψϚ� �Ͼ�a�������*� տ7�I�[��ϖߨߺ� ���߁���&�8�J� \��߀������s� ������k�4�F�X�j� |�������������� 0BT��	s ������� �>Pbt�)�������SCR�E?ǝ�u1sc�u2�3$33$43$53$6�3$73$83!#TAT~�� ֓+Ek��USER /,$k�s5#�$3�$4�$5*�$6�$7�$8�!s��NDO_CFG �X����s�PD�v!�)�N�one��� _IN_FO 1Y+EZ0Ԑ0%�u?�Hc? �?�?�?�?�?�?O�? 4OOXOjOMO�O�O�O��O��G1OFFSEOT \��^1�O ���_'_9_K_x_ o_�_�_�_�__�_o �_o>o5oGotoko}o@�o�[ן�m�o�o
�o|#�HUFRAM7���6D1RTO?L_ABRTGB3�_rENBhYxGR�P 1]�ӑCz  A��s�q1 ������(�:��[v��U�x1w{MSOK  �uZ1����[vNDq%R9�%�AXIS_6_�T��*�JR_EV�Ngp��6�22�^�K
 h1�UEVgp!td�:\event_�user\Џ+�C�70� 0Fe�#�S�P)�.�spot�weld`�!CA6��f�x���d!�o ?���2�ݗ���!�� e���E�W�Я{����� ��ï<��`���S� ����̿w������� 8����n�ϒϤ�Oπa��υ��ϩϻ� �W�RK 2_�)q8��b�t� Pߙ߫� �����߼�����;� M�(�q��^���� �������%� �6�[��m��$VARS__CONFI0`�K� FP��t�C7CRG2c�J�O�����DA��BeHJ�pC�J��*(?�: �$���MR�r2i�K�l�0	q���@�1: SC130EF2 *�� �e��X��ș��50�1<A@C�N�� �� �!NsIv�8�,0b� B���� �Z�:/�;/ &/_/J/�/n/�/�// �/�/�/�/%?�I?[?.��TCC��j�z@Ѝ98���j ��GF��
�k�K �%�UF12 Au�to �0 e s�et �R�� �h"u� 
�1em��~3456789'012I�A� ��0�����H�������fX�:��3�Q�.:$@8�@9� ~(:�o=L�@m���y���%I��O��j����%� ��O��1��_%W [B-hOzO�O�O�_�O �H�_�__%_'_9_K_ ]_o_�_no�_�_�o�_ �_�oo#o5oGo~�1�SELEC넙�����qVIA_WO�:�l���p��,�		��`�o�G��P ǫp�iXqSIONTMOU�� ��u��m��:��<t�1� FR:\�s\�DATA̟�0��� UD1:\ ��LOG�   �%��EX0�'� B@ ���s�D�iPen�dant 249� .design?.local;�[����= �� � n6  ����Ɯp��t#`φ	?  =����~� 
 MC�vTRAINZ��2��dO�p�����m�}��sOn�; (1[���
9������ џ���=�+�E�O��a�s�����z�ISS?TAT o�9y�� =-2997.�6665: wa�s less t�han acce�ptable v�alue: -1O00.0)���$80_SIDE_B4��g;IS_GE�sp6�;����
rpj |��\�HOMIN�p_q�E�����rHqq�aC$B�m�\�JMPERR {2r�;
  �o �����e���.�_�R� d�vψϚϬ������`���Dc�W�RE�p�s�|�LEXg�tܐ��@1-eP�VM�PHASE  ���j!r�OFF�SET_ENB��uOyP2�tu�KF��|���<�cB`A�1�`� ?s#33���1cA���cE��|��x���H�x��A����M� �j ��5�y��x<��t�9I�?��i� �����Ö0��Õ���[�{�3��1��� �E��҅�&��Z� �w?�1����Ⱦ��{� 1�������!S���# ��~������ �+ OAsh� ������
/ 9K]R/�'/�/ �/�/�/�]/�/5/*? <?k/]?�/i?�?�?�/ �?�/�??OC?U?�? EOSOeO{O�?�O�?�? 	O�O-O�O�O+_=_O_ y_�O	_{_�O�_�__ 	os_o?o9o�_xo�_ �o�_�o�_oKo�o�o�'5w[�TD_F�ILTE�yo�3 �f�t����o� �������'� 9�Ɓf�x����������ҏ����W�SH�IFTMENU [1z�<�%� f�1�D�j���z���ٟ �������W�.��@���d�v�ï��	�LIVE/SNA�P��vsfli�v��կ�b�I�ON ��U���menu����r����3�$���{b���M�O��|n��zY�W�AITDINEND  ��Kᷲ�sOK����OUT�r�S,���TIML���W�G�y�π��+�|�J�|�i���R�ELE������TM��˳���_AC�T���u���_DA�TA }b�v�%�  RIPPER_OPEN���`��RDIS1�-���$XS��~b������J���Z�XVR���;�$ZA�BC_GRP 1U����`,�h2��n�ZIP���F��sc�o������z�MPCF_G 1��� 0�o'���?�ك���`p��� 	�8�/�<�T�  �8U��?��;�\�����7iq����غ�����\���D��z�?��C2���5f��	����jv�
��e��&|��x�����������"��0������?{�^p|�f���b ����ݗ边�D#B���
�� � �
 .X�����:.@5��ৰ�����_CYLINuDfq��� Јf ,(  */�.-�c/W/>/{/b- ��/�/�./�/g/ ???R?�/v?�?�? �/�?Y???�?�?O�?`m?NO`O�?�2���x� ���O�o���O�_\�O8_�g��RQA��SPHE_RE 2��̲? �_O�_�_�_�_0OC_ o0o�?To�_�_�oqo �o�oo�o�o=oOo, �oP7I��o��l�9�ZZ�� ǳ�